// HwJSoC.v

// Generated using ACDS version 13.1 162 at 2020.06.26.19:30:19

`timescale 1 ps / 1 ps
module HwJSoC (
		input  wire        clk_clk,                      //                   clk.clk
		input  wire        reset_reset_n,                //                 reset.reset_n
		output wire        pll_c2_clk,                   //                pll_c2.clk
		output wire [7:0]  led_out_export,               //               led_out.export
		output wire [12:0] sdram_bus_addr,               //             sdram_bus.addr
		output wire [1:0]  sdram_bus_ba,                 //                      .ba
		output wire        sdram_bus_cas_n,              //                      .cas_n
		output wire        sdram_bus_cke,                //                      .cke
		output wire        sdram_bus_cs_n,               //                      .cs_n
		inout  wire [31:0] sdram_bus_dq,                 //                      .dq
		output wire [3:0]  sdram_bus_dqm,                //                      .dqm
		output wire        sdram_bus_ras_n,              //                      .ras_n
		output wire        sdram_bus_we_n,               //                      .we_n
		output wire        pll_c1_conduit_export,        //        pll_c1_conduit.export
		output wire        pll_locked_conduit_export,    //    pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export, // pll_phasedone_conduit.export
		input  wire        pll_areset_conduit_export     //    pll_areset_conduit.export
	);

	wire         pll_c0_clk;                                             // PLL:c0 -> [SDRAM_controller:clk, cpu_A:clk, cpu_B:clk, cpu_C:clk, cpu_D:clk, cpu_E:clk, cpu_F:clk, fifo_AB_0:wrclock, fifo_AB_1:wrclock, fifo_AB_2:wrclock, fifo_AD:wrclock, fifo_AE:wrclock, fifo_AF:wrclock, fifo_BC:wrclock, fifo_CD:wrclock, fifo_DE:wrclock, fifo_EF:wrclock, highTimer_A:clk, highTimer_B:clk, highTimer_C:clk, highTimer_D:clk, highTimer_E:clk, highTimer_F:clk, irq_mapper:clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_mapper_003:clk, irq_mapper_004:clk, irq_mapper_005:clk, jtag_A:clk, jtag_B:clk, jtag_C:clk, jtag_D:clk, jtag_E:clk, jtag_F:clk, led_out:clk, mm_interconnect_0:PLL_c0_clk, rst_controller:clk, rst_controller_002:clk, rst_controller_003:clk, rst_controller_004:clk, rst_controller_005:clk, rst_controller_006:clk, rst_controller_007:clk, rst_controller_008:clk, rst_controller_009:clk, rst_controller_010:clk, rst_controller_011:clk, rst_controller_012:clk, rst_controller_013:clk, rst_controller_014:clk, rst_controller_015:clk, sysid_A:clock, sysid_B:clock, sysid_C:clock, sysid_D:clock, sysid_E:clock, sysid_F:clock, timer_A:clk, timer_B:clk, timer_C:clk, timer_D:clk, timer_E:clk, timer_F:clk]
	wire         mm_interconnect_0_cpu_b_jtag_debug_module_waitrequest;  // cpu_B:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_B_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_b_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_B_jtag_debug_module_writedata -> cpu_B:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_b_jtag_debug_module_address;      // mm_interconnect_0:cpu_B_jtag_debug_module_address -> cpu_B:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_b_jtag_debug_module_write;        // mm_interconnect_0:cpu_B_jtag_debug_module_write -> cpu_B:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_b_jtag_debug_module_read;         // mm_interconnect_0:cpu_B_jtag_debug_module_read -> cpu_B:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_b_jtag_debug_module_readdata;     // cpu_B:jtag_debug_module_readdata -> mm_interconnect_0:cpu_B_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_b_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_B_jtag_debug_module_debugaccess -> cpu_B:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_b_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_B_jtag_debug_module_byteenable -> cpu_B:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_timer_d_s1_writedata;                 // mm_interconnect_0:timer_D_s1_writedata -> timer_D:writedata
	wire   [2:0] mm_interconnect_0_timer_d_s1_address;                   // mm_interconnect_0:timer_D_s1_address -> timer_D:address
	wire         mm_interconnect_0_timer_d_s1_chipselect;                // mm_interconnect_0:timer_D_s1_chipselect -> timer_D:chipselect
	wire         mm_interconnect_0_timer_d_s1_write;                     // mm_interconnect_0:timer_D_s1_write -> timer_D:write_n
	wire  [15:0] mm_interconnect_0_timer_d_s1_readdata;                  // timer_D:readdata -> mm_interconnect_0:timer_D_s1_readdata
	wire  [15:0] mm_interconnect_0_hightimer_c_s1_writedata;             // mm_interconnect_0:highTimer_C_s1_writedata -> highTimer_C:writedata
	wire   [2:0] mm_interconnect_0_hightimer_c_s1_address;               // mm_interconnect_0:highTimer_C_s1_address -> highTimer_C:address
	wire         mm_interconnect_0_hightimer_c_s1_chipselect;            // mm_interconnect_0:highTimer_C_s1_chipselect -> highTimer_C:chipselect
	wire         mm_interconnect_0_hightimer_c_s1_write;                 // mm_interconnect_0:highTimer_C_s1_write -> highTimer_C:write_n
	wire  [15:0] mm_interconnect_0_hightimer_c_s1_readdata;              // highTimer_C:readdata -> mm_interconnect_0:highTimer_C_s1_readdata
	wire  [31:0] mm_interconnect_0_fifo_ab_1_in_csr_writedata;           // mm_interconnect_0:fifo_AB_1_in_csr_writedata -> fifo_AB_1:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ab_1_in_csr_address;             // mm_interconnect_0:fifo_AB_1_in_csr_address -> fifo_AB_1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ab_1_in_csr_write;               // mm_interconnect_0:fifo_AB_1_in_csr_write -> fifo_AB_1:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ab_1_in_csr_read;                // mm_interconnect_0:fifo_AB_1_in_csr_read -> fifo_AB_1:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_1_in_csr_readdata;            // fifo_AB_1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AB_1_in_csr_readdata
	wire         mm_interconnect_0_jtag_e_avalon_jtag_slave_waitrequest; // jtag_E:av_waitrequest -> mm_interconnect_0:jtag_E_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_e_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_E_avalon_jtag_slave_writedata -> jtag_E:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_e_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_E_avalon_jtag_slave_address -> jtag_E:av_address
	wire         mm_interconnect_0_jtag_e_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_E_avalon_jtag_slave_chipselect -> jtag_E:av_chipselect
	wire         mm_interconnect_0_jtag_e_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_E_avalon_jtag_slave_write -> jtag_E:av_write_n
	wire         mm_interconnect_0_jtag_e_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_E_avalon_jtag_slave_read -> jtag_E:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_e_avalon_jtag_slave_readdata;    // jtag_E:av_readdata -> mm_interconnect_0:jtag_E_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo_de_in_csr_writedata;             // mm_interconnect_0:fifo_DE_in_csr_writedata -> fifo_DE:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_de_in_csr_address;               // mm_interconnect_0:fifo_DE_in_csr_address -> fifo_DE:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_de_in_csr_write;                 // mm_interconnect_0:fifo_DE_in_csr_write -> fifo_DE:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_de_in_csr_read;                  // mm_interconnect_0:fifo_DE_in_csr_read -> fifo_DE:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_de_in_csr_readdata;              // fifo_DE:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_DE_in_csr_readdata
	wire  [31:0] mm_interconnect_0_fifo_ef_in_csr_writedata;             // mm_interconnect_0:fifo_EF_in_csr_writedata -> fifo_EF:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ef_in_csr_address;               // mm_interconnect_0:fifo_EF_in_csr_address -> fifo_EF:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ef_in_csr_write;                 // mm_interconnect_0:fifo_EF_in_csr_write -> fifo_EF:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ef_in_csr_read;                  // mm_interconnect_0:fifo_EF_in_csr_read -> fifo_EF:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ef_in_csr_readdata;              // fifo_EF:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_EF_in_csr_readdata
	wire         cpu_d_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_D_instruction_master_waitrequest -> cpu_D:i_waitrequest
	wire  [27:0] cpu_d_instruction_master_address;                       // cpu_D:i_address -> mm_interconnect_0:cpu_D_instruction_master_address
	wire         cpu_d_instruction_master_read;                          // cpu_D:i_read -> mm_interconnect_0:cpu_D_instruction_master_read
	wire  [31:0] cpu_d_instruction_master_readdata;                      // mm_interconnect_0:cpu_D_instruction_master_readdata -> cpu_D:i_readdata
	wire         cpu_d_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_D_instruction_master_readdatavalid -> cpu_D:i_readdatavalid
	wire         cpu_d_data_master_waitrequest;                          // mm_interconnect_0:cpu_D_data_master_waitrequest -> cpu_D:d_waitrequest
	wire  [31:0] cpu_d_data_master_writedata;                            // cpu_D:d_writedata -> mm_interconnect_0:cpu_D_data_master_writedata
	wire  [27:0] cpu_d_data_master_address;                              // cpu_D:d_address -> mm_interconnect_0:cpu_D_data_master_address
	wire         cpu_d_data_master_write;                                // cpu_D:d_write -> mm_interconnect_0:cpu_D_data_master_write
	wire         cpu_d_data_master_read;                                 // cpu_D:d_read -> mm_interconnect_0:cpu_D_data_master_read
	wire  [31:0] cpu_d_data_master_readdata;                             // mm_interconnect_0:cpu_D_data_master_readdata -> cpu_D:d_readdata
	wire         cpu_d_data_master_debugaccess;                          // cpu_D:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_D_data_master_debugaccess
	wire   [3:0] cpu_d_data_master_byteenable;                           // cpu_D:d_byteenable -> mm_interconnect_0:cpu_D_data_master_byteenable
	wire         cpu_c_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_C_instruction_master_waitrequest -> cpu_C:i_waitrequest
	wire  [27:0] cpu_c_instruction_master_address;                       // cpu_C:i_address -> mm_interconnect_0:cpu_C_instruction_master_address
	wire         cpu_c_instruction_master_read;                          // cpu_C:i_read -> mm_interconnect_0:cpu_C_instruction_master_read
	wire  [31:0] cpu_c_instruction_master_readdata;                      // mm_interconnect_0:cpu_C_instruction_master_readdata -> cpu_C:i_readdata
	wire         cpu_c_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_C_instruction_master_readdatavalid -> cpu_C:i_readdatavalid
	wire         cpu_f_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_F_instruction_master_waitrequest -> cpu_F:i_waitrequest
	wire  [27:0] cpu_f_instruction_master_address;                       // cpu_F:i_address -> mm_interconnect_0:cpu_F_instruction_master_address
	wire         cpu_f_instruction_master_read;                          // cpu_F:i_read -> mm_interconnect_0:cpu_F_instruction_master_read
	wire  [31:0] cpu_f_instruction_master_readdata;                      // mm_interconnect_0:cpu_F_instruction_master_readdata -> cpu_F:i_readdata
	wire         cpu_f_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_F_instruction_master_readdatavalid -> cpu_F:i_readdatavalid
	wire         cpu_e_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_E_instruction_master_waitrequest -> cpu_E:i_waitrequest
	wire  [27:0] cpu_e_instruction_master_address;                       // cpu_E:i_address -> mm_interconnect_0:cpu_E_instruction_master_address
	wire         cpu_e_instruction_master_read;                          // cpu_E:i_read -> mm_interconnect_0:cpu_E_instruction_master_read
	wire  [31:0] cpu_e_instruction_master_readdata;                      // mm_interconnect_0:cpu_E_instruction_master_readdata -> cpu_E:i_readdata
	wire         cpu_e_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_E_instruction_master_readdatavalid -> cpu_E:i_readdatavalid
	wire         mm_interconnect_0_fifo_ab_1_in_waitrequest;             // fifo_AB_1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AB_1_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ab_1_in_writedata;               // mm_interconnect_0:fifo_AB_1_in_writedata -> fifo_AB_1:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ab_1_in_write;                   // mm_interconnect_0:fifo_AB_1_in_write -> fifo_AB_1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_ab_0_in_csr_writedata;           // mm_interconnect_0:fifo_AB_0_in_csr_writedata -> fifo_AB_0:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ab_0_in_csr_address;             // mm_interconnect_0:fifo_AB_0_in_csr_address -> fifo_AB_0:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ab_0_in_csr_write;               // mm_interconnect_0:fifo_AB_0_in_csr_write -> fifo_AB_0:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ab_0_in_csr_read;                // mm_interconnect_0:fifo_AB_0_in_csr_read -> fifo_AB_0:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_0_in_csr_readdata;            // fifo_AB_0:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AB_0_in_csr_readdata
	wire         mm_interconnect_0_fifo_ae_in_waitrequest;               // fifo_AE:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AE_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ae_in_writedata;                 // mm_interconnect_0:fifo_AE_in_writedata -> fifo_AE:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ae_in_write;                     // mm_interconnect_0:fifo_AE_in_write -> fifo_AE:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_ad_out_waitrequest;              // fifo_AD:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AD_out_waitrequest
	wire         mm_interconnect_0_fifo_ad_out_read;                     // mm_interconnect_0:fifo_AD_out_read -> fifo_AD:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ad_out_readdata;                 // fifo_AD:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AD_out_readdata
	wire         mm_interconnect_0_fifo_ad_in_waitrequest;               // fifo_AD:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AD_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ad_in_writedata;                 // mm_interconnect_0:fifo_AD_in_writedata -> fifo_AD:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ad_in_write;                     // mm_interconnect_0:fifo_AD_in_write -> fifo_AD:avalonmm_write_slave_write
	wire   [0:0] mm_interconnect_0_sysid_a_control_slave_address;        // mm_interconnect_0:sysid_A_control_slave_address -> sysid_A:address
	wire  [31:0] mm_interconnect_0_sysid_a_control_slave_readdata;       // sysid_A:readdata -> mm_interconnect_0:sysid_A_control_slave_readdata
	wire  [15:0] mm_interconnect_0_hightimer_f_s1_writedata;             // mm_interconnect_0:highTimer_F_s1_writedata -> highTimer_F:writedata
	wire   [2:0] mm_interconnect_0_hightimer_f_s1_address;               // mm_interconnect_0:highTimer_F_s1_address -> highTimer_F:address
	wire         mm_interconnect_0_hightimer_f_s1_chipselect;            // mm_interconnect_0:highTimer_F_s1_chipselect -> highTimer_F:chipselect
	wire         mm_interconnect_0_hightimer_f_s1_write;                 // mm_interconnect_0:highTimer_F_s1_write -> highTimer_F:write_n
	wire  [15:0] mm_interconnect_0_hightimer_f_s1_readdata;              // highTimer_F:readdata -> mm_interconnect_0:highTimer_F_s1_readdata
	wire         mm_interconnect_0_fifo_cd_in_waitrequest;               // fifo_CD:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_CD_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_cd_in_writedata;                 // mm_interconnect_0:fifo_CD_in_writedata -> fifo_CD:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_cd_in_write;                     // mm_interconnect_0:fifo_CD_in_write -> fifo_CD:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_ef_out_waitrequest;              // fifo_EF:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_EF_out_waitrequest
	wire         mm_interconnect_0_fifo_ef_out_read;                     // mm_interconnect_0:fifo_EF_out_read -> fifo_EF:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ef_out_readdata;                 // fifo_EF:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_EF_out_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;      // SDRAM_controller:za_waitrequest -> mm_interconnect_0:SDRAM_controller_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;        // mm_interconnect_0:SDRAM_controller_s1_writedata -> SDRAM_controller:az_data
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;          // mm_interconnect_0:SDRAM_controller_s1_address -> SDRAM_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;       // mm_interconnect_0:SDRAM_controller_s1_chipselect -> SDRAM_controller:az_cs
	wire         mm_interconnect_0_sdram_controller_s1_write;            // mm_interconnect_0:SDRAM_controller_s1_write -> SDRAM_controller:az_wr_n
	wire         mm_interconnect_0_sdram_controller_s1_read;             // mm_interconnect_0:SDRAM_controller_s1_read -> SDRAM_controller:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;         // SDRAM_controller:za_data -> mm_interconnect_0:SDRAM_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;    // SDRAM_controller:za_valid -> mm_interconnect_0:SDRAM_controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;       // mm_interconnect_0:SDRAM_controller_s1_byteenable -> SDRAM_controller:az_be_n
	wire         mm_interconnect_0_fifo_af_in_waitrequest;               // fifo_AF:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AF_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_af_in_writedata;                 // mm_interconnect_0:fifo_AF_in_writedata -> fifo_AF:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_af_in_write;                     // mm_interconnect_0:fifo_AF_in_write -> fifo_AF:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_ab_0_out_waitrequest;            // fifo_AB_0:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AB_0_out_waitrequest
	wire         mm_interconnect_0_fifo_ab_0_out_read;                   // mm_interconnect_0:fifo_AB_0_out_read -> fifo_AB_0:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_0_out_readdata;               // fifo_AB_0:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AB_0_out_readdata
	wire         mm_interconnect_0_fifo_ab_2_in_waitrequest;             // fifo_AB_2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AB_2_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ab_2_in_writedata;               // mm_interconnect_0:fifo_AB_2_in_writedata -> fifo_AB_2:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ab_2_in_write;                   // mm_interconnect_0:fifo_AB_2_in_write -> fifo_AB_2:avalonmm_write_slave_write
	wire         cpu_e_data_master_waitrequest;                          // mm_interconnect_0:cpu_E_data_master_waitrequest -> cpu_E:d_waitrequest
	wire  [31:0] cpu_e_data_master_writedata;                            // cpu_E:d_writedata -> mm_interconnect_0:cpu_E_data_master_writedata
	wire  [27:0] cpu_e_data_master_address;                              // cpu_E:d_address -> mm_interconnect_0:cpu_E_data_master_address
	wire         cpu_e_data_master_write;                                // cpu_E:d_write -> mm_interconnect_0:cpu_E_data_master_write
	wire         cpu_e_data_master_read;                                 // cpu_E:d_read -> mm_interconnect_0:cpu_E_data_master_read
	wire  [31:0] cpu_e_data_master_readdata;                             // mm_interconnect_0:cpu_E_data_master_readdata -> cpu_E:d_readdata
	wire         cpu_e_data_master_debugaccess;                          // cpu_E:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_E_data_master_debugaccess
	wire   [3:0] cpu_e_data_master_byteenable;                           // cpu_E:d_byteenable -> mm_interconnect_0:cpu_E_data_master_byteenable
	wire         cpu_b_data_master_waitrequest;                          // mm_interconnect_0:cpu_B_data_master_waitrequest -> cpu_B:d_waitrequest
	wire  [31:0] cpu_b_data_master_writedata;                            // cpu_B:d_writedata -> mm_interconnect_0:cpu_B_data_master_writedata
	wire  [27:0] cpu_b_data_master_address;                              // cpu_B:d_address -> mm_interconnect_0:cpu_B_data_master_address
	wire         cpu_b_data_master_write;                                // cpu_B:d_write -> mm_interconnect_0:cpu_B_data_master_write
	wire         cpu_b_data_master_read;                                 // cpu_B:d_read -> mm_interconnect_0:cpu_B_data_master_read
	wire  [31:0] cpu_b_data_master_readdata;                             // mm_interconnect_0:cpu_B_data_master_readdata -> cpu_B:d_readdata
	wire         cpu_b_data_master_debugaccess;                          // cpu_B:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_B_data_master_debugaccess
	wire   [3:0] cpu_b_data_master_byteenable;                           // cpu_B:d_byteenable -> mm_interconnect_0:cpu_B_data_master_byteenable
	wire  [31:0] mm_interconnect_0_fifo_ad_in_csr_writedata;             // mm_interconnect_0:fifo_AD_in_csr_writedata -> fifo_AD:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ad_in_csr_address;               // mm_interconnect_0:fifo_AD_in_csr_address -> fifo_AD:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ad_in_csr_write;                 // mm_interconnect_0:fifo_AD_in_csr_write -> fifo_AD:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ad_in_csr_read;                  // mm_interconnect_0:fifo_AD_in_csr_read -> fifo_AD:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ad_in_csr_readdata;              // fifo_AD:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AD_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer_e_s1_writedata;                 // mm_interconnect_0:timer_E_s1_writedata -> timer_E:writedata
	wire   [2:0] mm_interconnect_0_timer_e_s1_address;                   // mm_interconnect_0:timer_E_s1_address -> timer_E:address
	wire         mm_interconnect_0_timer_e_s1_chipselect;                // mm_interconnect_0:timer_E_s1_chipselect -> timer_E:chipselect
	wire         mm_interconnect_0_timer_e_s1_write;                     // mm_interconnect_0:timer_E_s1_write -> timer_E:write_n
	wire  [15:0] mm_interconnect_0_timer_e_s1_readdata;                  // timer_E:readdata -> mm_interconnect_0:timer_E_s1_readdata
	wire         mm_interconnect_0_fifo_ef_in_waitrequest;               // fifo_EF:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_EF_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ef_in_writedata;                 // mm_interconnect_0:fifo_EF_in_writedata -> fifo_EF:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ef_in_write;                     // mm_interconnect_0:fifo_EF_in_write -> fifo_EF:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_ae_in_csr_writedata;             // mm_interconnect_0:fifo_AE_in_csr_writedata -> fifo_AE:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ae_in_csr_address;               // mm_interconnect_0:fifo_AE_in_csr_address -> fifo_AE:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ae_in_csr_write;                 // mm_interconnect_0:fifo_AE_in_csr_write -> fifo_AE:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ae_in_csr_read;                  // mm_interconnect_0:fifo_AE_in_csr_read -> fifo_AE:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ae_in_csr_readdata;              // fifo_AE:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AE_in_csr_readdata
	wire         mm_interconnect_0_fifo_bc_out_waitrequest;              // fifo_BC:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_BC_out_waitrequest
	wire         mm_interconnect_0_fifo_bc_out_read;                     // mm_interconnect_0:fifo_BC_out_read -> fifo_BC:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_bc_out_readdata;                 // fifo_BC:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_BC_out_readdata
	wire  [15:0] mm_interconnect_0_timer_c_s1_writedata;                 // mm_interconnect_0:timer_C_s1_writedata -> timer_C:writedata
	wire   [2:0] mm_interconnect_0_timer_c_s1_address;                   // mm_interconnect_0:timer_C_s1_address -> timer_C:address
	wire         mm_interconnect_0_timer_c_s1_chipselect;                // mm_interconnect_0:timer_C_s1_chipselect -> timer_C:chipselect
	wire         mm_interconnect_0_timer_c_s1_write;                     // mm_interconnect_0:timer_C_s1_write -> timer_C:write_n
	wire  [15:0] mm_interconnect_0_timer_c_s1_readdata;                  // timer_C:readdata -> mm_interconnect_0:timer_C_s1_readdata
	wire  [15:0] mm_interconnect_0_hightimer_b_s1_writedata;             // mm_interconnect_0:highTimer_B_s1_writedata -> highTimer_B:writedata
	wire   [2:0] mm_interconnect_0_hightimer_b_s1_address;               // mm_interconnect_0:highTimer_B_s1_address -> highTimer_B:address
	wire         mm_interconnect_0_hightimer_b_s1_chipselect;            // mm_interconnect_0:highTimer_B_s1_chipselect -> highTimer_B:chipselect
	wire         mm_interconnect_0_hightimer_b_s1_write;                 // mm_interconnect_0:highTimer_B_s1_write -> highTimer_B:write_n
	wire  [15:0] mm_interconnect_0_hightimer_b_s1_readdata;              // highTimer_B:readdata -> mm_interconnect_0:highTimer_B_s1_readdata
	wire         cpu_f_data_master_waitrequest;                          // mm_interconnect_0:cpu_F_data_master_waitrequest -> cpu_F:d_waitrequest
	wire  [31:0] cpu_f_data_master_writedata;                            // cpu_F:d_writedata -> mm_interconnect_0:cpu_F_data_master_writedata
	wire  [27:0] cpu_f_data_master_address;                              // cpu_F:d_address -> mm_interconnect_0:cpu_F_data_master_address
	wire         cpu_f_data_master_write;                                // cpu_F:d_write -> mm_interconnect_0:cpu_F_data_master_write
	wire         cpu_f_data_master_read;                                 // cpu_F:d_read -> mm_interconnect_0:cpu_F_data_master_read
	wire  [31:0] cpu_f_data_master_readdata;                             // mm_interconnect_0:cpu_F_data_master_readdata -> cpu_F:d_readdata
	wire         cpu_f_data_master_debugaccess;                          // cpu_F:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_F_data_master_debugaccess
	wire   [3:0] cpu_f_data_master_byteenable;                           // cpu_F:d_byteenable -> mm_interconnect_0:cpu_F_data_master_byteenable
	wire         cpu_a_data_master_waitrequest;                          // mm_interconnect_0:cpu_A_data_master_waitrequest -> cpu_A:d_waitrequest
	wire  [31:0] cpu_a_data_master_writedata;                            // cpu_A:d_writedata -> mm_interconnect_0:cpu_A_data_master_writedata
	wire  [27:0] cpu_a_data_master_address;                              // cpu_A:d_address -> mm_interconnect_0:cpu_A_data_master_address
	wire         cpu_a_data_master_write;                                // cpu_A:d_write -> mm_interconnect_0:cpu_A_data_master_write
	wire         cpu_a_data_master_read;                                 // cpu_A:d_read -> mm_interconnect_0:cpu_A_data_master_read
	wire  [31:0] cpu_a_data_master_readdata;                             // mm_interconnect_0:cpu_A_data_master_readdata -> cpu_A:d_readdata
	wire         cpu_a_data_master_debugaccess;                          // cpu_A:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_A_data_master_debugaccess
	wire   [3:0] cpu_a_data_master_byteenable;                           // cpu_A:d_byteenable -> mm_interconnect_0:cpu_A_data_master_byteenable
	wire         mm_interconnect_0_jtag_d_avalon_jtag_slave_waitrequest; // jtag_D:av_waitrequest -> mm_interconnect_0:jtag_D_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_d_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_D_avalon_jtag_slave_writedata -> jtag_D:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_d_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_D_avalon_jtag_slave_address -> jtag_D:av_address
	wire         mm_interconnect_0_jtag_d_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_D_avalon_jtag_slave_chipselect -> jtag_D:av_chipselect
	wire         mm_interconnect_0_jtag_d_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_D_avalon_jtag_slave_write -> jtag_D:av_write_n
	wire         mm_interconnect_0_jtag_d_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_D_avalon_jtag_slave_read -> jtag_D:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_d_avalon_jtag_slave_readdata;    // jtag_D:av_readdata -> mm_interconnect_0:jtag_D_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_fifo_ab_2_out_waitrequest;            // fifo_AB_2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AB_2_out_waitrequest
	wire         mm_interconnect_0_fifo_ab_2_out_read;                   // mm_interconnect_0:fifo_AB_2_out_read -> fifo_AB_2:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_2_out_readdata;               // fifo_AB_2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AB_2_out_readdata
	wire         mm_interconnect_0_cpu_d_jtag_debug_module_waitrequest;  // cpu_D:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_D_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_d_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_D_jtag_debug_module_writedata -> cpu_D:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_d_jtag_debug_module_address;      // mm_interconnect_0:cpu_D_jtag_debug_module_address -> cpu_D:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_d_jtag_debug_module_write;        // mm_interconnect_0:cpu_D_jtag_debug_module_write -> cpu_D:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_d_jtag_debug_module_read;         // mm_interconnect_0:cpu_D_jtag_debug_module_read -> cpu_D:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_d_jtag_debug_module_readdata;     // cpu_D:jtag_debug_module_readdata -> mm_interconnect_0:cpu_D_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_d_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_D_jtag_debug_module_debugaccess -> cpu_D:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_d_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_D_jtag_debug_module_byteenable -> cpu_D:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_fifo_cd_in_csr_writedata;             // mm_interconnect_0:fifo_CD_in_csr_writedata -> fifo_CD:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_cd_in_csr_address;               // mm_interconnect_0:fifo_CD_in_csr_address -> fifo_CD:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_cd_in_csr_write;                 // mm_interconnect_0:fifo_CD_in_csr_write -> fifo_CD:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_cd_in_csr_read;                  // mm_interconnect_0:fifo_CD_in_csr_read -> fifo_CD:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_cd_in_csr_readdata;              // fifo_CD:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_CD_in_csr_readdata
	wire   [0:0] mm_interconnect_0_sysid_d_control_slave_address;        // mm_interconnect_0:sysid_D_control_slave_address -> sysid_D:address
	wire  [31:0] mm_interconnect_0_sysid_d_control_slave_readdata;       // sysid_D:readdata -> mm_interconnect_0:sysid_D_control_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_b_s1_writedata;                 // mm_interconnect_0:timer_B_s1_writedata -> timer_B:writedata
	wire   [2:0] mm_interconnect_0_timer_b_s1_address;                   // mm_interconnect_0:timer_B_s1_address -> timer_B:address
	wire         mm_interconnect_0_timer_b_s1_chipselect;                // mm_interconnect_0:timer_B_s1_chipselect -> timer_B:chipselect
	wire         mm_interconnect_0_timer_b_s1_write;                     // mm_interconnect_0:timer_B_s1_write -> timer_B:write_n
	wire  [15:0] mm_interconnect_0_timer_b_s1_readdata;                  // timer_B:readdata -> mm_interconnect_0:timer_B_s1_readdata
	wire         mm_interconnect_0_fifo_bc_in_waitrequest;               // fifo_BC:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_BC_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_bc_in_writedata;                 // mm_interconnect_0:fifo_BC_in_writedata -> fifo_BC:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_bc_in_write;                     // mm_interconnect_0:fifo_BC_in_write -> fifo_BC:avalonmm_write_slave_write
	wire   [0:0] mm_interconnect_0_sysid_c_control_slave_address;        // mm_interconnect_0:sysid_C_control_slave_address -> sysid_C:address
	wire  [31:0] mm_interconnect_0_sysid_c_control_slave_readdata;       // sysid_C:readdata -> mm_interconnect_0:sysid_C_control_slave_readdata
	wire         mm_interconnect_0_cpu_f_jtag_debug_module_waitrequest;  // cpu_F:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_F_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_f_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_F_jtag_debug_module_writedata -> cpu_F:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_f_jtag_debug_module_address;      // mm_interconnect_0:cpu_F_jtag_debug_module_address -> cpu_F:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_f_jtag_debug_module_write;        // mm_interconnect_0:cpu_F_jtag_debug_module_write -> cpu_F:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_f_jtag_debug_module_read;         // mm_interconnect_0:cpu_F_jtag_debug_module_read -> cpu_F:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_f_jtag_debug_module_readdata;     // cpu_F:jtag_debug_module_readdata -> mm_interconnect_0:cpu_F_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_f_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_F_jtag_debug_module_debugaccess -> cpu_F:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_f_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_F_jtag_debug_module_byteenable -> cpu_F:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo_cd_out_waitrequest;              // fifo_CD:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_CD_out_waitrequest
	wire         mm_interconnect_0_fifo_cd_out_read;                     // mm_interconnect_0:fifo_CD_out_read -> fifo_CD:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_cd_out_readdata;                 // fifo_CD:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_CD_out_readdata
	wire         mm_interconnect_0_fifo_ab_0_in_waitrequest;             // fifo_AB_0:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_AB_0_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_ab_0_in_writedata;               // mm_interconnect_0:fifo_AB_0_in_writedata -> fifo_AB_0:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_ab_0_in_write;                   // mm_interconnect_0:fifo_AB_0_in_write -> fifo_AB_0:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_ab_2_in_csr_writedata;           // mm_interconnect_0:fifo_AB_2_in_csr_writedata -> fifo_AB_2:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_ab_2_in_csr_address;             // mm_interconnect_0:fifo_AB_2_in_csr_address -> fifo_AB_2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_ab_2_in_csr_write;               // mm_interconnect_0:fifo_AB_2_in_csr_write -> fifo_AB_2:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_ab_2_in_csr_read;                // mm_interconnect_0:fifo_AB_2_in_csr_read -> fifo_AB_2:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_2_in_csr_readdata;            // fifo_AB_2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AB_2_in_csr_readdata
	wire         mm_interconnect_0_jtag_c_avalon_jtag_slave_waitrequest; // jtag_C:av_waitrequest -> mm_interconnect_0:jtag_C_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_c_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_C_avalon_jtag_slave_writedata -> jtag_C:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_c_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_C_avalon_jtag_slave_address -> jtag_C:av_address
	wire         mm_interconnect_0_jtag_c_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_C_avalon_jtag_slave_chipselect -> jtag_C:av_chipselect
	wire         mm_interconnect_0_jtag_c_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_C_avalon_jtag_slave_write -> jtag_C:av_write_n
	wire         mm_interconnect_0_jtag_c_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_C_avalon_jtag_slave_read -> jtag_C:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_c_avalon_jtag_slave_readdata;    // jtag_C:av_readdata -> mm_interconnect_0:jtag_C_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_b_avalon_jtag_slave_waitrequest; // jtag_B:av_waitrequest -> mm_interconnect_0:jtag_B_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_b_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_B_avalon_jtag_slave_writedata -> jtag_B:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_b_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_B_avalon_jtag_slave_address -> jtag_B:av_address
	wire         mm_interconnect_0_jtag_b_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_B_avalon_jtag_slave_chipselect -> jtag_B:av_chipselect
	wire         mm_interconnect_0_jtag_b_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_B_avalon_jtag_slave_write -> jtag_B:av_write_n
	wire         mm_interconnect_0_jtag_b_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_B_avalon_jtag_slave_read -> jtag_B:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_b_avalon_jtag_slave_readdata;    // jtag_B:av_readdata -> mm_interconnect_0:jtag_B_avalon_jtag_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_b_control_slave_address;        // mm_interconnect_0:sysid_B_control_slave_address -> sysid_B:address
	wire  [31:0] mm_interconnect_0_sysid_b_control_slave_readdata;       // sysid_B:readdata -> mm_interconnect_0:sysid_B_control_slave_readdata
	wire  [15:0] mm_interconnect_0_hightimer_a_s1_writedata;             // mm_interconnect_0:highTimer_A_s1_writedata -> highTimer_A:writedata
	wire   [2:0] mm_interconnect_0_hightimer_a_s1_address;               // mm_interconnect_0:highTimer_A_s1_address -> highTimer_A:address
	wire         mm_interconnect_0_hightimer_a_s1_chipselect;            // mm_interconnect_0:highTimer_A_s1_chipselect -> highTimer_A:chipselect
	wire         mm_interconnect_0_hightimer_a_s1_write;                 // mm_interconnect_0:highTimer_A_s1_write -> highTimer_A:write_n
	wire  [15:0] mm_interconnect_0_hightimer_a_s1_readdata;              // highTimer_A:readdata -> mm_interconnect_0:highTimer_A_s1_readdata
	wire         mm_interconnect_0_fifo_de_out_waitrequest;              // fifo_DE:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_DE_out_waitrequest
	wire         mm_interconnect_0_fifo_de_out_read;                     // mm_interconnect_0:fifo_DE_out_read -> fifo_DE:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_de_out_readdata;                 // fifo_DE:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_DE_out_readdata
	wire  [15:0] mm_interconnect_0_hightimer_d_s1_writedata;             // mm_interconnect_0:highTimer_D_s1_writedata -> highTimer_D:writedata
	wire   [2:0] mm_interconnect_0_hightimer_d_s1_address;               // mm_interconnect_0:highTimer_D_s1_address -> highTimer_D:address
	wire         mm_interconnect_0_hightimer_d_s1_chipselect;            // mm_interconnect_0:highTimer_D_s1_chipselect -> highTimer_D:chipselect
	wire         mm_interconnect_0_hightimer_d_s1_write;                 // mm_interconnect_0:highTimer_D_s1_write -> highTimer_D:write_n
	wire  [15:0] mm_interconnect_0_hightimer_d_s1_readdata;              // highTimer_D:readdata -> mm_interconnect_0:highTimer_D_s1_readdata
	wire  [15:0] mm_interconnect_0_hightimer_e_s1_writedata;             // mm_interconnect_0:highTimer_E_s1_writedata -> highTimer_E:writedata
	wire   [2:0] mm_interconnect_0_hightimer_e_s1_address;               // mm_interconnect_0:highTimer_E_s1_address -> highTimer_E:address
	wire         mm_interconnect_0_hightimer_e_s1_chipselect;            // mm_interconnect_0:highTimer_E_s1_chipselect -> highTimer_E:chipselect
	wire         mm_interconnect_0_hightimer_e_s1_write;                 // mm_interconnect_0:highTimer_E_s1_write -> highTimer_E:write_n
	wire  [15:0] mm_interconnect_0_hightimer_e_s1_readdata;              // highTimer_E:readdata -> mm_interconnect_0:highTimer_E_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_e_control_slave_address;        // mm_interconnect_0:sysid_E_control_slave_address -> sysid_E:address
	wire  [31:0] mm_interconnect_0_sysid_e_control_slave_readdata;       // sysid_E:readdata -> mm_interconnect_0:sysid_E_control_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_a_s1_writedata;                 // mm_interconnect_0:timer_A_s1_writedata -> timer_A:writedata
	wire   [2:0] mm_interconnect_0_timer_a_s1_address;                   // mm_interconnect_0:timer_A_s1_address -> timer_A:address
	wire         mm_interconnect_0_timer_a_s1_chipselect;                // mm_interconnect_0:timer_A_s1_chipselect -> timer_A:chipselect
	wire         mm_interconnect_0_timer_a_s1_write;                     // mm_interconnect_0:timer_A_s1_write -> timer_A:write_n
	wire  [15:0] mm_interconnect_0_timer_a_s1_readdata;                  // timer_A:readdata -> mm_interconnect_0:timer_A_s1_readdata
	wire         mm_interconnect_0_fifo_ae_out_waitrequest;              // fifo_AE:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AE_out_waitrequest
	wire         mm_interconnect_0_fifo_ae_out_read;                     // mm_interconnect_0:fifo_AE_out_read -> fifo_AE:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ae_out_readdata;                 // fifo_AE:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AE_out_readdata
	wire         mm_interconnect_0_cpu_a_jtag_debug_module_waitrequest;  // cpu_A:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_A_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_a_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_A_jtag_debug_module_writedata -> cpu_A:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_a_jtag_debug_module_address;      // mm_interconnect_0:cpu_A_jtag_debug_module_address -> cpu_A:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_a_jtag_debug_module_write;        // mm_interconnect_0:cpu_A_jtag_debug_module_write -> cpu_A:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_a_jtag_debug_module_read;         // mm_interconnect_0:cpu_A_jtag_debug_module_read -> cpu_A:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_a_jtag_debug_module_readdata;     // cpu_A:jtag_debug_module_readdata -> mm_interconnect_0:cpu_A_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_a_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_A_jtag_debug_module_debugaccess -> cpu_A:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_a_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_A_jtag_debug_module_byteenable -> cpu_A:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo_af_out_waitrequest;              // fifo_AF:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AF_out_waitrequest
	wire         mm_interconnect_0_fifo_af_out_read;                     // mm_interconnect_0:fifo_AF_out_read -> fifo_AF:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_af_out_readdata;                 // fifo_AF:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AF_out_readdata
	wire         mm_interconnect_0_fifo_de_in_waitrequest;               // fifo_DE:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_DE_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_de_in_writedata;                 // mm_interconnect_0:fifo_DE_in_writedata -> fifo_DE:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_de_in_write;                     // mm_interconnect_0:fifo_DE_in_write -> fifo_DE:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_ab_1_out_waitrequest;            // fifo_AB_1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_AB_1_out_waitrequest
	wire         mm_interconnect_0_fifo_ab_1_out_read;                   // mm_interconnect_0:fifo_AB_1_out_read -> fifo_AB_1:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_ab_1_out_readdata;               // fifo_AB_1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_AB_1_out_readdata
	wire         cpu_b_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_B_instruction_master_waitrequest -> cpu_B:i_waitrequest
	wire  [27:0] cpu_b_instruction_master_address;                       // cpu_B:i_address -> mm_interconnect_0:cpu_B_instruction_master_address
	wire         cpu_b_instruction_master_read;                          // cpu_B:i_read -> mm_interconnect_0:cpu_B_instruction_master_read
	wire  [31:0] cpu_b_instruction_master_readdata;                      // mm_interconnect_0:cpu_B_instruction_master_readdata -> cpu_B:i_readdata
	wire         cpu_b_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_B_instruction_master_readdatavalid -> cpu_B:i_readdatavalid
	wire         mm_interconnect_0_jtag_f_avalon_jtag_slave_waitrequest; // jtag_F:av_waitrequest -> mm_interconnect_0:jtag_F_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_f_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_F_avalon_jtag_slave_writedata -> jtag_F:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_f_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_F_avalon_jtag_slave_address -> jtag_F:av_address
	wire         mm_interconnect_0_jtag_f_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_F_avalon_jtag_slave_chipselect -> jtag_F:av_chipselect
	wire         mm_interconnect_0_jtag_f_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_F_avalon_jtag_slave_write -> jtag_F:av_write_n
	wire         mm_interconnect_0_jtag_f_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_F_avalon_jtag_slave_read -> jtag_F:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_f_avalon_jtag_slave_readdata;    // jtag_F:av_readdata -> mm_interconnect_0:jtag_F_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo_af_in_csr_writedata;             // mm_interconnect_0:fifo_AF_in_csr_writedata -> fifo_AF:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_af_in_csr_address;               // mm_interconnect_0:fifo_AF_in_csr_address -> fifo_AF:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_af_in_csr_write;                 // mm_interconnect_0:fifo_AF_in_csr_write -> fifo_AF:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_af_in_csr_read;                  // mm_interconnect_0:fifo_AF_in_csr_read -> fifo_AF:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_af_in_csr_readdata;              // fifo_AF:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_AF_in_csr_readdata
	wire  [31:0] mm_interconnect_0_fifo_bc_in_csr_writedata;             // mm_interconnect_0:fifo_BC_in_csr_writedata -> fifo_BC:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_bc_in_csr_address;               // mm_interconnect_0:fifo_BC_in_csr_address -> fifo_BC:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_bc_in_csr_write;                 // mm_interconnect_0:fifo_BC_in_csr_write -> fifo_BC:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_bc_in_csr_read;                  // mm_interconnect_0:fifo_BC_in_csr_read -> fifo_BC:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_bc_in_csr_readdata;              // fifo_BC:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_BC_in_csr_readdata
	wire   [0:0] mm_interconnect_0_sysid_f_control_slave_address;        // mm_interconnect_0:sysid_F_control_slave_address -> sysid_F:address
	wire  [31:0] mm_interconnect_0_sysid_f_control_slave_readdata;       // sysid_F:readdata -> mm_interconnect_0:sysid_F_control_slave_readdata
	wire  [31:0] mm_interconnect_0_led_out_s1_writedata;                 // mm_interconnect_0:led_out_s1_writedata -> led_out:writedata
	wire   [1:0] mm_interconnect_0_led_out_s1_address;                   // mm_interconnect_0:led_out_s1_address -> led_out:address
	wire         mm_interconnect_0_led_out_s1_chipselect;                // mm_interconnect_0:led_out_s1_chipselect -> led_out:chipselect
	wire         mm_interconnect_0_led_out_s1_write;                     // mm_interconnect_0:led_out_s1_write -> led_out:write_n
	wire  [31:0] mm_interconnect_0_led_out_s1_readdata;                  // led_out:readdata -> mm_interconnect_0:led_out_s1_readdata
	wire         mm_interconnect_0_cpu_c_jtag_debug_module_waitrequest;  // cpu_C:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_C_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_c_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_C_jtag_debug_module_writedata -> cpu_C:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_c_jtag_debug_module_address;      // mm_interconnect_0:cpu_C_jtag_debug_module_address -> cpu_C:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_c_jtag_debug_module_write;        // mm_interconnect_0:cpu_C_jtag_debug_module_write -> cpu_C:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_c_jtag_debug_module_read;         // mm_interconnect_0:cpu_C_jtag_debug_module_read -> cpu_C:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_c_jtag_debug_module_readdata;     // cpu_C:jtag_debug_module_readdata -> mm_interconnect_0:cpu_C_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_c_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_C_jtag_debug_module_debugaccess -> cpu_C:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_c_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_C_jtag_debug_module_byteenable -> cpu_C:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_e_jtag_debug_module_waitrequest;  // cpu_E:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_E_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_e_jtag_debug_module_writedata;    // mm_interconnect_0:cpu_E_jtag_debug_module_writedata -> cpu_E:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_e_jtag_debug_module_address;      // mm_interconnect_0:cpu_E_jtag_debug_module_address -> cpu_E:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_e_jtag_debug_module_write;        // mm_interconnect_0:cpu_E_jtag_debug_module_write -> cpu_E:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_e_jtag_debug_module_read;         // mm_interconnect_0:cpu_E_jtag_debug_module_read -> cpu_E:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_e_jtag_debug_module_readdata;     // cpu_E:jtag_debug_module_readdata -> mm_interconnect_0:cpu_E_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_e_jtag_debug_module_debugaccess;  // mm_interconnect_0:cpu_E_jtag_debug_module_debugaccess -> cpu_E:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_e_jtag_debug_module_byteenable;   // mm_interconnect_0:cpu_E_jtag_debug_module_byteenable -> cpu_E:jtag_debug_module_byteenable
	wire         cpu_a_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_A_instruction_master_waitrequest -> cpu_A:i_waitrequest
	wire  [27:0] cpu_a_instruction_master_address;                       // cpu_A:i_address -> mm_interconnect_0:cpu_A_instruction_master_address
	wire         cpu_a_instruction_master_read;                          // cpu_A:i_read -> mm_interconnect_0:cpu_A_instruction_master_read
	wire  [31:0] cpu_a_instruction_master_readdata;                      // mm_interconnect_0:cpu_A_instruction_master_readdata -> cpu_A:i_readdata
	wire         cpu_a_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_A_instruction_master_readdatavalid -> cpu_A:i_readdatavalid
	wire         mm_interconnect_0_jtag_a_avalon_jtag_slave_waitrequest; // jtag_A:av_waitrequest -> mm_interconnect_0:jtag_A_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_a_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_A_avalon_jtag_slave_writedata -> jtag_A:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_a_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_A_avalon_jtag_slave_address -> jtag_A:av_address
	wire         mm_interconnect_0_jtag_a_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_A_avalon_jtag_slave_chipselect -> jtag_A:av_chipselect
	wire         mm_interconnect_0_jtag_a_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_A_avalon_jtag_slave_write -> jtag_A:av_write_n
	wire         mm_interconnect_0_jtag_a_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_A_avalon_jtag_slave_read -> jtag_A:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_a_avalon_jtag_slave_readdata;    // jtag_A:av_readdata -> mm_interconnect_0:jtag_A_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_f_s1_writedata;                 // mm_interconnect_0:timer_F_s1_writedata -> timer_F:writedata
	wire   [2:0] mm_interconnect_0_timer_f_s1_address;                   // mm_interconnect_0:timer_F_s1_address -> timer_F:address
	wire         mm_interconnect_0_timer_f_s1_chipselect;                // mm_interconnect_0:timer_F_s1_chipselect -> timer_F:chipselect
	wire         mm_interconnect_0_timer_f_s1_write;                     // mm_interconnect_0:timer_F_s1_write -> timer_F:write_n
	wire  [15:0] mm_interconnect_0_timer_f_s1_readdata;                  // timer_F:readdata -> mm_interconnect_0:timer_F_s1_readdata
	wire         cpu_c_data_master_waitrequest;                          // mm_interconnect_0:cpu_C_data_master_waitrequest -> cpu_C:d_waitrequest
	wire  [31:0] cpu_c_data_master_writedata;                            // cpu_C:d_writedata -> mm_interconnect_0:cpu_C_data_master_writedata
	wire  [27:0] cpu_c_data_master_address;                              // cpu_C:d_address -> mm_interconnect_0:cpu_C_data_master_address
	wire         cpu_c_data_master_write;                                // cpu_C:d_write -> mm_interconnect_0:cpu_C_data_master_write
	wire         cpu_c_data_master_read;                                 // cpu_C:d_read -> mm_interconnect_0:cpu_C_data_master_read
	wire  [31:0] cpu_c_data_master_readdata;                             // mm_interconnect_0:cpu_C_data_master_readdata -> cpu_C:d_readdata
	wire         cpu_c_data_master_debugaccess;                          // cpu_C:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_C_data_master_debugaccess
	wire   [3:0] cpu_c_data_master_byteenable;                           // cpu_C:d_byteenable -> mm_interconnect_0:cpu_C_data_master_byteenable
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;              // mm_interconnect_0:PLL_pll_slave_writedata -> PLL:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                // mm_interconnect_0:PLL_pll_slave_address -> PLL:address
	wire         mm_interconnect_0_pll_pll_slave_write;                  // mm_interconnect_0:PLL_pll_slave_write -> PLL:write
	wire         mm_interconnect_0_pll_pll_slave_read;                   // mm_interconnect_0:PLL_pll_slave_read -> PLL:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;               // PLL:readdata -> mm_interconnect_0:PLL_pll_slave_readdata
	wire         irq_mapper_receiver0_irq;                               // timer_A:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                               // jtag_A:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                               // highTimer_A:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                               // fifo_AB_0:wrclk_control_slave_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                               // fifo_AB_2:wrclk_control_slave_irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                               // fifo_AB_1:wrclk_control_slave_irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver7_irq;                               // fifo_AF:wrclk_control_slave_irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                               // fifo_AE:wrclk_control_slave_irq -> irq_mapper:receiver8_irq
	wire  [31:0] cpu_a_d_irq_irq;                                        // irq_mapper:sender_irq -> cpu_A:d_irq
	wire         irq_mapper_001_receiver0_irq;                           // highTimer_B:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                           // timer_B:irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver2_irq;                           // jtag_B:av_irq -> irq_mapper_001:receiver2_irq
	wire         irq_mapper_001_receiver3_irq;                           // fifo_BC:wrclk_control_slave_irq -> irq_mapper_001:receiver3_irq
	wire  [31:0] cpu_b_d_irq_irq;                                        // irq_mapper_001:sender_irq -> cpu_B:d_irq
	wire         irq_mapper_002_receiver0_irq;                           // timer_C:irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                           // highTimer_C:irq -> irq_mapper_002:receiver1_irq
	wire         irq_mapper_002_receiver2_irq;                           // jtag_C:av_irq -> irq_mapper_002:receiver2_irq
	wire         irq_mapper_002_receiver3_irq;                           // fifo_CD:wrclk_control_slave_irq -> irq_mapper_002:receiver3_irq
	wire  [31:0] cpu_c_d_irq_irq;                                        // irq_mapper_002:sender_irq -> cpu_C:d_irq
	wire         irq_mapper_003_receiver0_irq;                           // timer_D:irq -> irq_mapper_003:receiver0_irq
	wire         irq_mapper_003_receiver1_irq;                           // highTimer_D:irq -> irq_mapper_003:receiver1_irq
	wire         irq_mapper_003_receiver2_irq;                           // jtag_D:av_irq -> irq_mapper_003:receiver2_irq
	wire         irq_mapper_003_receiver3_irq;                           // fifo_DE:wrclk_control_slave_irq -> irq_mapper_003:receiver3_irq
	wire  [31:0] cpu_d_d_irq_irq;                                        // irq_mapper_003:sender_irq -> cpu_D:d_irq
	wire         irq_mapper_004_receiver0_irq;                           // timer_E:irq -> irq_mapper_004:receiver0_irq
	wire         irq_mapper_004_receiver1_irq;                           // highTimer_E:irq -> irq_mapper_004:receiver1_irq
	wire         irq_mapper_004_receiver2_irq;                           // jtag_E:av_irq -> irq_mapper_004:receiver2_irq
	wire         irq_mapper_004_receiver3_irq;                           // fifo_EF:wrclk_control_slave_irq -> irq_mapper_004:receiver3_irq
	wire  [31:0] cpu_e_d_irq_irq;                                        // irq_mapper_004:sender_irq -> cpu_E:d_irq
	wire         irq_mapper_005_receiver0_irq;                           // timer_F:irq -> irq_mapper_005:receiver0_irq
	wire         irq_mapper_005_receiver1_irq;                           // highTimer_F:irq -> irq_mapper_005:receiver1_irq
	wire         irq_mapper_005_receiver2_irq;                           // jtag_F:av_irq -> irq_mapper_005:receiver2_irq
	wire  [31:0] cpu_f_d_irq_irq;                                        // irq_mapper_005:sender_irq -> cpu_F:d_irq
	wire         irq_mapper_receiver6_irq;                               // fifo_AD:wrclk_control_slave_irq -> [irq_mapper:receiver6_irq, irq_mapper_003:receiver4_irq]
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [SDRAM_controller:reset_n, led_out:reset_n, mm_interconnect_0:SDRAM_controller_reset_reset_bridge_in_reset_reset]
	wire         cpu_a_jtag_debug_module_reset_reset;                    // cpu_A:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_002:reset_in0, rst_controller_003:reset_in1, rst_controller_009:reset_in1, rst_controller_010:reset_in1, rst_controller_011:reset_in1]
	wire         cpu_c_jtag_debug_module_reset_reset;                    // cpu_C:jtag_debug_module_resetrequest -> [rst_controller:reset_in2, rst_controller_005:reset_in0, rst_controller_012:reset_in2, rst_controller_013:reset_in1]
	wire         cpu_d_jtag_debug_module_reset_reset;                    // cpu_D:jtag_debug_module_resetrequest -> [rst_controller:reset_in3, rst_controller_006:reset_in0, rst_controller_009:reset_in2, rst_controller_013:reset_in2, rst_controller_014:reset_in1]
	wire         cpu_b_jtag_debug_module_reset_reset;                    // cpu_B:jtag_debug_module_resetrequest -> [rst_controller:reset_in4, rst_controller_003:reset_in2, rst_controller_004:reset_in1, rst_controller_012:reset_in1]
	wire         cpu_e_jtag_debug_module_reset_reset;                    // cpu_E:jtag_debug_module_resetrequest -> [rst_controller:reset_in5, rst_controller_007:reset_in0, rst_controller_010:reset_in2, rst_controller_014:reset_in2, rst_controller_015:reset_in0]
	wire         cpu_f_jtag_debug_module_reset_reset;                    // cpu_F:jtag_debug_module_resetrequest -> [rst_controller:reset_in6, rst_controller_008:reset_in0, rst_controller_011:reset_in2, rst_controller_015:reset_in2]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [PLL:reset, mm_interconnect_0:PLL_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                     // rst_controller_002:reset_out -> [cpu_A:reset_n, highTimer_A:reset_n, irq_mapper:reset, jtag_A:rst_n, mm_interconnect_0:cpu_A_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid_A:reset_n, timer_A:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                 // rst_controller_002:reset_req -> [cpu_A:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                     // rst_controller_003:reset_out -> [fifo_AB_0:reset_n, fifo_AB_1:reset_n, fifo_AB_2:reset_n, mm_interconnect_0:fifo_AB_0_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                     // rst_controller_004:reset_out -> [cpu_B:reset_n, highTimer_B:reset_n, irq_mapper_001:reset, jtag_B:rst_n, mm_interconnect_0:cpu_B_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset, sysid_B:reset_n, timer_B:reset_n]
	wire         rst_controller_004_reset_out_reset_req;                 // rst_controller_004:reset_req -> [cpu_B:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_005_reset_out_reset;                     // rst_controller_005:reset_out -> [cpu_C:reset_n, highTimer_C:reset_n, irq_mapper_002:reset, jtag_C:rst_n, mm_interconnect_0:cpu_C_reset_n_reset_bridge_in_reset_reset, rst_translator_002:in_reset, sysid_C:reset_n, timer_C:reset_n]
	wire         rst_controller_005_reset_out_reset_req;                 // rst_controller_005:reset_req -> [cpu_C:reset_req, rst_translator_002:reset_req_in]
	wire         rst_controller_006_reset_out_reset;                     // rst_controller_006:reset_out -> [cpu_D:reset_n, highTimer_D:reset_n, irq_mapper_003:reset, jtag_D:rst_n, mm_interconnect_0:cpu_D_reset_n_reset_bridge_in_reset_reset, rst_translator_003:in_reset, sysid_D:reset_n, timer_D:reset_n]
	wire         rst_controller_006_reset_out_reset_req;                 // rst_controller_006:reset_req -> [cpu_D:reset_req, rst_translator_003:reset_req_in]
	wire         rst_controller_007_reset_out_reset;                     // rst_controller_007:reset_out -> [cpu_E:reset_n, highTimer_E:reset_n, irq_mapper_004:reset, jtag_E:rst_n, mm_interconnect_0:cpu_E_reset_n_reset_bridge_in_reset_reset, rst_translator_004:in_reset, sysid_E:reset_n, timer_E:reset_n]
	wire         rst_controller_007_reset_out_reset_req;                 // rst_controller_007:reset_req -> [cpu_E:reset_req, rst_translator_004:reset_req_in]
	wire         rst_controller_008_reset_out_reset;                     // rst_controller_008:reset_out -> [cpu_F:reset_n, highTimer_F:reset_n, irq_mapper_005:reset, jtag_F:rst_n, mm_interconnect_0:cpu_F_reset_n_reset_bridge_in_reset_reset, rst_translator_005:in_reset, sysid_F:reset_n, timer_F:reset_n]
	wire         rst_controller_008_reset_out_reset_req;                 // rst_controller_008:reset_req -> [cpu_F:reset_req, rst_translator_005:reset_req_in]
	wire         rst_controller_009_reset_out_reset;                     // rst_controller_009:reset_out -> [fifo_AD:reset_n, mm_interconnect_0:fifo_AD_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_010_reset_out_reset;                     // rst_controller_010:reset_out -> [fifo_AE:reset_n, mm_interconnect_0:fifo_AE_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_011_reset_out_reset;                     // rst_controller_011:reset_out -> [fifo_AF:reset_n, mm_interconnect_0:fifo_AF_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_012_reset_out_reset;                     // rst_controller_012:reset_out -> [fifo_BC:reset_n, mm_interconnect_0:fifo_BC_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_013_reset_out_reset;                     // rst_controller_013:reset_out -> [fifo_CD:reset_n, mm_interconnect_0:fifo_CD_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_014_reset_out_reset;                     // rst_controller_014:reset_out -> [fifo_DE:reset_n, mm_interconnect_0:fifo_DE_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_015_reset_out_reset;                     // rst_controller_015:reset_out -> [fifo_EF:reset_n, mm_interconnect_0:fifo_EF_reset_in_reset_bridge_in_reset_reset]

	HwJSoC_SDRAM_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_bus_addr),                                      //  wire.export
		.zs_ba          (sdram_bus_ba),                                        //      .export
		.zs_cas_n       (sdram_bus_cas_n),                                     //      .export
		.zs_cke         (sdram_bus_cke),                                       //      .export
		.zs_cs_n        (sdram_bus_cs_n),                                      //      .export
		.zs_dq          (sdram_bus_dq),                                        //      .export
		.zs_dqm         (sdram_bus_dqm),                                       //      .export
		.zs_ras_n       (sdram_bus_ras_n),                                     //      .export
		.zs_we_n        (sdram_bus_we_n)                                       //      .export
	);

	HwJSoC_PLL pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c2        (pll_c2_clk),                                //                    c2.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.c1        (pll_c1_conduit_export),                     //            c1_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	HwJSoC_led_out led_out (
		.clk        (pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_out_s1_readdata),   //                    .readdata
		.out_port   (led_out_export)                           // external_connection.export
	);

	HwJSoC_timer_A timer_a (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_a_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_a_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_a_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_a_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_a_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_a (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_a_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_a_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_a (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_a_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_a_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_a_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_a_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_a_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_a_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_a_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                //               irq.irq
	);

	HwJSoC_cpu_A cpu_a (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_a_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_a_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_a_data_master_read),                                //                          .read
		.d_readdata                            (cpu_a_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_a_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_a_data_master_write),                               //                          .write
		.d_writedata                           (cpu_a_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_a_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_a_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_a_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_a_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_a_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_a_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_a_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_a_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_a_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_a_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_a_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_a_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_a_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_a_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_a_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_a_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_highTimer_A hightimer_a (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_a_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_a_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_a_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_a_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_a_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                     //   irq.irq
	);

	HwJSoC_fifo_AB_0 fifo_ab_0 (
		.wrclock                          (pll_c0_clk),                                   //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ab_0_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ab_0_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ab_0_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ab_0_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ab_0_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ab_0_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ab_0_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ab_0_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ab_0_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ab_0_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ab_0_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver3_irq)                      //   in_irq.irq
	);

	HwJSoC_timer_A timer_b (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_b_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_b_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_b_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_b_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_b_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver1_irq)             //   irq.irq
	);

	HwJSoC_highTimer_A hightimer_b (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_b_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_b_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_b_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_b_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_b_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_b (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_b_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_b_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_b (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_b_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_b_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_b_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_b_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_b_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_b_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_b_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver2_irq)                            //               irq.irq
	);

	HwJSoC_cpu_B cpu_b (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_004_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_004_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_b_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_b_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_b_data_master_read),                                //                          .read
		.d_readdata                            (cpu_b_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_b_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_b_data_master_write),                               //                          .write
		.d_writedata                           (cpu_b_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_b_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_b_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_b_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_b_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_b_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_b_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_b_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_b_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_b_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_b_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_b_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_b_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_b_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_b_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_b_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_b_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_timer_A timer_c (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_c_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_c_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_c_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_c_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_c_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)             //   irq.irq
	);

	HwJSoC_highTimer_A hightimer_c (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_c_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_c_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_c_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_c_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_c_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver1_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_c (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_c_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_c_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_c (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_005_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_c_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_c_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_c_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_c_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_c_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_c_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_c_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver2_irq)                            //               irq.irq
	);

	HwJSoC_cpu_C cpu_c (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_005_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_005_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_c_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_c_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_c_data_master_read),                                //                          .read
		.d_readdata                            (cpu_c_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_c_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_c_data_master_write),                               //                          .write
		.d_writedata                           (cpu_c_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_c_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_c_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_c_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_c_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_c_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_c_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_c_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_c_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_c_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_c_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_c_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_c_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_c_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_c_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_c_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_c_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_timer_A timer_d (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_d_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_d_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_d_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_d_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_d_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver0_irq)             //   irq.irq
	);

	HwJSoC_highTimer_A hightimer_d (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_d_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_d_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_d_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_d_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_d_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver1_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_d (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_006_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_d_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_d_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_d (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_006_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_d_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_d_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_d_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_d_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_d_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_d_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_d_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver2_irq)                            //               irq.irq
	);

	HwJSoC_cpu_D cpu_d (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_006_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_006_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_d_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_d_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_d_data_master_read),                                //                          .read
		.d_readdata                            (cpu_d_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_d_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_d_data_master_write),                               //                          .write
		.d_writedata                           (cpu_d_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_d_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_d_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_d_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_d_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_d_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_d_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_d_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_d_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_d_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_d_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_d_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_d_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_d_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_d_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_d_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_timer_A timer_e (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_007_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_e_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_e_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_e_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_e_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_e_s1_write),     //      .write_n
		.irq        (irq_mapper_004_receiver0_irq)             //   irq.irq
	);

	HwJSoC_highTimer_A hightimer_e (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_007_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_e_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_e_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_e_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_e_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_e_s1_write),     //      .write_n
		.irq        (irq_mapper_004_receiver1_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_e (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_007_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_e_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_e_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_e (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_007_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_e_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_e_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_e_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_e_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_e_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_e_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_e_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_004_receiver2_irq)                            //               irq.irq
	);

	HwJSoC_cpu_E cpu_e (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_007_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_007_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_e_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_e_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_e_data_master_read),                                //                          .read
		.d_readdata                            (cpu_e_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_e_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_e_data_master_write),                               //                          .write
		.d_writedata                           (cpu_e_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_e_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_e_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_e_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_e_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_e_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_e_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_e_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_e_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_e_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_e_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_e_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_e_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_e_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_e_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_e_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_e_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_timer_A timer_f (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_008_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_f_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_f_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_f_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_f_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_f_s1_write),     //      .write_n
		.irq        (irq_mapper_005_receiver0_irq)             //   irq.irq
	);

	HwJSoC_highTimer_A hightimer_f (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_008_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_hightimer_f_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hightimer_f_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hightimer_f_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hightimer_f_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hightimer_f_s1_write),     //      .write_n
		.irq        (irq_mapper_005_receiver1_irq)                 //   irq.irq
	);

	HwJSoC_sysid_A sysid_f (
		.clock    (pll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_008_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_f_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_f_control_slave_address)   //              .address
	);

	HwJSoC_jtag_A jtag_f (
		.clk            (pll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_008_reset_out_reset),                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_f_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_f_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_f_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_f_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_f_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_f_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_f_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_005_receiver2_irq)                            //               irq.irq
	);

	HwJSoC_cpu_F cpu_f (
		.clk                                   (pll_c0_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_008_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_008_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_f_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_f_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_f_data_master_read),                                //                          .read
		.d_readdata                            (cpu_f_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_f_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_f_data_master_write),                               //                          .write
		.d_writedata                           (cpu_f_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_f_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_f_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_f_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_f_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_f_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_f_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_f_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_f_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_f_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_f_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_f_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_f_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_f_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_f_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_f_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_f_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	HwJSoC_fifo_AB_0 fifo_ab_1 (
		.wrclock                          (pll_c0_clk),                                   //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ab_1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ab_1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ab_1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ab_1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ab_1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ab_1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ab_1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ab_1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ab_1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ab_1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ab_1_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver5_irq)                      //   in_irq.irq
	);

	HwJSoC_fifo_AB_0 fifo_ab_2 (
		.wrclock                          (pll_c0_clk),                                   //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ab_2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ab_2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ab_2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ab_2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ab_2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ab_2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ab_2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ab_2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ab_2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ab_2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ab_2_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver4_irq)                      //   in_irq.irq
	);

	HwJSoC_fifo_AD fifo_ad (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_009_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ad_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ad_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ad_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ad_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ad_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ad_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ad_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ad_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ad_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ad_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ad_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver6_irq)                    //   in_irq.irq
	);

	HwJSoC_fifo_AD fifo_ae (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_010_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ae_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ae_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ae_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ae_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ae_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ae_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ae_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ae_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ae_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ae_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ae_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver8_irq)                    //   in_irq.irq
	);

	HwJSoC_fifo_AD fifo_af (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_011_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_af_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_af_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_af_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_af_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_af_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_af_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_af_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_af_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_af_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_af_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_af_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver7_irq)                    //   in_irq.irq
	);

	HwJSoC_fifo_BC fifo_bc (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_012_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_bc_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_bc_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_bc_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_bc_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_bc_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_bc_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_bc_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_bc_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_bc_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_bc_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_bc_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_001_receiver3_irq)                //   in_irq.irq
	);

	HwJSoC_fifo_BC fifo_cd (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_013_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_cd_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_cd_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_cd_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_cd_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_cd_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_cd_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_cd_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_cd_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_cd_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_cd_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_cd_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_002_receiver3_irq)                //   in_irq.irq
	);

	HwJSoC_fifo_BC fifo_de (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_014_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_de_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_de_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_de_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_de_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_de_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_de_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_de_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_de_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_de_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_de_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_de_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_003_receiver3_irq)                //   in_irq.irq
	);

	HwJSoC_fifo_EF fifo_ef (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_015_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_ef_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_ef_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_ef_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_ef_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_ef_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_ef_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_ef_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_ef_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_ef_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_ef_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_ef_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_004_receiver3_irq)                //   in_irq.irq
	);

	HwJSoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clk_clk),                                                //                                       clock_clk.clk
		.PLL_c0_clk                                            (pll_c0_clk),                                             //                                          PLL_c0.clk
		.cpu_A_reset_n_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                     //             cpu_A_reset_n_reset_bridge_in_reset.reset
		.cpu_B_reset_n_reset_bridge_in_reset_reset             (rst_controller_004_reset_out_reset),                     //             cpu_B_reset_n_reset_bridge_in_reset.reset
		.cpu_C_reset_n_reset_bridge_in_reset_reset             (rst_controller_005_reset_out_reset),                     //             cpu_C_reset_n_reset_bridge_in_reset.reset
		.cpu_D_reset_n_reset_bridge_in_reset_reset             (rst_controller_006_reset_out_reset),                     //             cpu_D_reset_n_reset_bridge_in_reset.reset
		.cpu_E_reset_n_reset_bridge_in_reset_reset             (rst_controller_007_reset_out_reset),                     //             cpu_E_reset_n_reset_bridge_in_reset.reset
		.cpu_F_reset_n_reset_bridge_in_reset_reset             (rst_controller_008_reset_out_reset),                     //             cpu_F_reset_n_reset_bridge_in_reset.reset
		.fifo_AB_0_reset_in_reset_bridge_in_reset_reset        (rst_controller_003_reset_out_reset),                     //        fifo_AB_0_reset_in_reset_bridge_in_reset.reset
		.fifo_AD_reset_in_reset_bridge_in_reset_reset          (rst_controller_009_reset_out_reset),                     //          fifo_AD_reset_in_reset_bridge_in_reset.reset
		.fifo_AE_reset_in_reset_bridge_in_reset_reset          (rst_controller_010_reset_out_reset),                     //          fifo_AE_reset_in_reset_bridge_in_reset.reset
		.fifo_AF_reset_in_reset_bridge_in_reset_reset          (rst_controller_011_reset_out_reset),                     //          fifo_AF_reset_in_reset_bridge_in_reset.reset
		.fifo_BC_reset_in_reset_bridge_in_reset_reset          (rst_controller_012_reset_out_reset),                     //          fifo_BC_reset_in_reset_bridge_in_reset.reset
		.fifo_CD_reset_in_reset_bridge_in_reset_reset          (rst_controller_013_reset_out_reset),                     //          fifo_CD_reset_in_reset_bridge_in_reset.reset
		.fifo_DE_reset_in_reset_bridge_in_reset_reset          (rst_controller_014_reset_out_reset),                     //          fifo_DE_reset_in_reset_bridge_in_reset.reset
		.fifo_EF_reset_in_reset_bridge_in_reset_reset          (rst_controller_015_reset_out_reset),                     //          fifo_EF_reset_in_reset_bridge_in_reset.reset
		.PLL_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // PLL_inclk_interface_reset_reset_bridge_in_reset.reset
		.SDRAM_controller_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                         //    SDRAM_controller_reset_reset_bridge_in_reset.reset
		.cpu_A_data_master_address                             (cpu_a_data_master_address),                              //                               cpu_A_data_master.address
		.cpu_A_data_master_waitrequest                         (cpu_a_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_A_data_master_byteenable                          (cpu_a_data_master_byteenable),                           //                                                .byteenable
		.cpu_A_data_master_read                                (cpu_a_data_master_read),                                 //                                                .read
		.cpu_A_data_master_readdata                            (cpu_a_data_master_readdata),                             //                                                .readdata
		.cpu_A_data_master_write                               (cpu_a_data_master_write),                                //                                                .write
		.cpu_A_data_master_writedata                           (cpu_a_data_master_writedata),                            //                                                .writedata
		.cpu_A_data_master_debugaccess                         (cpu_a_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_A_instruction_master_address                      (cpu_a_instruction_master_address),                       //                        cpu_A_instruction_master.address
		.cpu_A_instruction_master_waitrequest                  (cpu_a_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_A_instruction_master_read                         (cpu_a_instruction_master_read),                          //                                                .read
		.cpu_A_instruction_master_readdata                     (cpu_a_instruction_master_readdata),                      //                                                .readdata
		.cpu_A_instruction_master_readdatavalid                (cpu_a_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_B_data_master_address                             (cpu_b_data_master_address),                              //                               cpu_B_data_master.address
		.cpu_B_data_master_waitrequest                         (cpu_b_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_B_data_master_byteenable                          (cpu_b_data_master_byteenable),                           //                                                .byteenable
		.cpu_B_data_master_read                                (cpu_b_data_master_read),                                 //                                                .read
		.cpu_B_data_master_readdata                            (cpu_b_data_master_readdata),                             //                                                .readdata
		.cpu_B_data_master_write                               (cpu_b_data_master_write),                                //                                                .write
		.cpu_B_data_master_writedata                           (cpu_b_data_master_writedata),                            //                                                .writedata
		.cpu_B_data_master_debugaccess                         (cpu_b_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_B_instruction_master_address                      (cpu_b_instruction_master_address),                       //                        cpu_B_instruction_master.address
		.cpu_B_instruction_master_waitrequest                  (cpu_b_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_B_instruction_master_read                         (cpu_b_instruction_master_read),                          //                                                .read
		.cpu_B_instruction_master_readdata                     (cpu_b_instruction_master_readdata),                      //                                                .readdata
		.cpu_B_instruction_master_readdatavalid                (cpu_b_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_C_data_master_address                             (cpu_c_data_master_address),                              //                               cpu_C_data_master.address
		.cpu_C_data_master_waitrequest                         (cpu_c_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_C_data_master_byteenable                          (cpu_c_data_master_byteenable),                           //                                                .byteenable
		.cpu_C_data_master_read                                (cpu_c_data_master_read),                                 //                                                .read
		.cpu_C_data_master_readdata                            (cpu_c_data_master_readdata),                             //                                                .readdata
		.cpu_C_data_master_write                               (cpu_c_data_master_write),                                //                                                .write
		.cpu_C_data_master_writedata                           (cpu_c_data_master_writedata),                            //                                                .writedata
		.cpu_C_data_master_debugaccess                         (cpu_c_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_C_instruction_master_address                      (cpu_c_instruction_master_address),                       //                        cpu_C_instruction_master.address
		.cpu_C_instruction_master_waitrequest                  (cpu_c_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_C_instruction_master_read                         (cpu_c_instruction_master_read),                          //                                                .read
		.cpu_C_instruction_master_readdata                     (cpu_c_instruction_master_readdata),                      //                                                .readdata
		.cpu_C_instruction_master_readdatavalid                (cpu_c_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_D_data_master_address                             (cpu_d_data_master_address),                              //                               cpu_D_data_master.address
		.cpu_D_data_master_waitrequest                         (cpu_d_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_D_data_master_byteenable                          (cpu_d_data_master_byteenable),                           //                                                .byteenable
		.cpu_D_data_master_read                                (cpu_d_data_master_read),                                 //                                                .read
		.cpu_D_data_master_readdata                            (cpu_d_data_master_readdata),                             //                                                .readdata
		.cpu_D_data_master_write                               (cpu_d_data_master_write),                                //                                                .write
		.cpu_D_data_master_writedata                           (cpu_d_data_master_writedata),                            //                                                .writedata
		.cpu_D_data_master_debugaccess                         (cpu_d_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_D_instruction_master_address                      (cpu_d_instruction_master_address),                       //                        cpu_D_instruction_master.address
		.cpu_D_instruction_master_waitrequest                  (cpu_d_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_D_instruction_master_read                         (cpu_d_instruction_master_read),                          //                                                .read
		.cpu_D_instruction_master_readdata                     (cpu_d_instruction_master_readdata),                      //                                                .readdata
		.cpu_D_instruction_master_readdatavalid                (cpu_d_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_E_data_master_address                             (cpu_e_data_master_address),                              //                               cpu_E_data_master.address
		.cpu_E_data_master_waitrequest                         (cpu_e_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_E_data_master_byteenable                          (cpu_e_data_master_byteenable),                           //                                                .byteenable
		.cpu_E_data_master_read                                (cpu_e_data_master_read),                                 //                                                .read
		.cpu_E_data_master_readdata                            (cpu_e_data_master_readdata),                             //                                                .readdata
		.cpu_E_data_master_write                               (cpu_e_data_master_write),                                //                                                .write
		.cpu_E_data_master_writedata                           (cpu_e_data_master_writedata),                            //                                                .writedata
		.cpu_E_data_master_debugaccess                         (cpu_e_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_E_instruction_master_address                      (cpu_e_instruction_master_address),                       //                        cpu_E_instruction_master.address
		.cpu_E_instruction_master_waitrequest                  (cpu_e_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_E_instruction_master_read                         (cpu_e_instruction_master_read),                          //                                                .read
		.cpu_E_instruction_master_readdata                     (cpu_e_instruction_master_readdata),                      //                                                .readdata
		.cpu_E_instruction_master_readdatavalid                (cpu_e_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_F_data_master_address                             (cpu_f_data_master_address),                              //                               cpu_F_data_master.address
		.cpu_F_data_master_waitrequest                         (cpu_f_data_master_waitrequest),                          //                                                .waitrequest
		.cpu_F_data_master_byteenable                          (cpu_f_data_master_byteenable),                           //                                                .byteenable
		.cpu_F_data_master_read                                (cpu_f_data_master_read),                                 //                                                .read
		.cpu_F_data_master_readdata                            (cpu_f_data_master_readdata),                             //                                                .readdata
		.cpu_F_data_master_write                               (cpu_f_data_master_write),                                //                                                .write
		.cpu_F_data_master_writedata                           (cpu_f_data_master_writedata),                            //                                                .writedata
		.cpu_F_data_master_debugaccess                         (cpu_f_data_master_debugaccess),                          //                                                .debugaccess
		.cpu_F_instruction_master_address                      (cpu_f_instruction_master_address),                       //                        cpu_F_instruction_master.address
		.cpu_F_instruction_master_waitrequest                  (cpu_f_instruction_master_waitrequest),                   //                                                .waitrequest
		.cpu_F_instruction_master_read                         (cpu_f_instruction_master_read),                          //                                                .read
		.cpu_F_instruction_master_readdata                     (cpu_f_instruction_master_readdata),                      //                                                .readdata
		.cpu_F_instruction_master_readdatavalid                (cpu_f_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.cpu_A_jtag_debug_module_address                       (mm_interconnect_0_cpu_a_jtag_debug_module_address),      //                         cpu_A_jtag_debug_module.address
		.cpu_A_jtag_debug_module_write                         (mm_interconnect_0_cpu_a_jtag_debug_module_write),        //                                                .write
		.cpu_A_jtag_debug_module_read                          (mm_interconnect_0_cpu_a_jtag_debug_module_read),         //                                                .read
		.cpu_A_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_a_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_A_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_a_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_A_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_a_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_A_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_a_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_A_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_a_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.cpu_B_jtag_debug_module_address                       (mm_interconnect_0_cpu_b_jtag_debug_module_address),      //                         cpu_B_jtag_debug_module.address
		.cpu_B_jtag_debug_module_write                         (mm_interconnect_0_cpu_b_jtag_debug_module_write),        //                                                .write
		.cpu_B_jtag_debug_module_read                          (mm_interconnect_0_cpu_b_jtag_debug_module_read),         //                                                .read
		.cpu_B_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_b_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_B_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_b_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_B_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_b_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_B_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_b_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_B_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_b_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.cpu_C_jtag_debug_module_address                       (mm_interconnect_0_cpu_c_jtag_debug_module_address),      //                         cpu_C_jtag_debug_module.address
		.cpu_C_jtag_debug_module_write                         (mm_interconnect_0_cpu_c_jtag_debug_module_write),        //                                                .write
		.cpu_C_jtag_debug_module_read                          (mm_interconnect_0_cpu_c_jtag_debug_module_read),         //                                                .read
		.cpu_C_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_c_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_C_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_c_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_C_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_c_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_C_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_c_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_C_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_c_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.cpu_D_jtag_debug_module_address                       (mm_interconnect_0_cpu_d_jtag_debug_module_address),      //                         cpu_D_jtag_debug_module.address
		.cpu_D_jtag_debug_module_write                         (mm_interconnect_0_cpu_d_jtag_debug_module_write),        //                                                .write
		.cpu_D_jtag_debug_module_read                          (mm_interconnect_0_cpu_d_jtag_debug_module_read),         //                                                .read
		.cpu_D_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_d_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_D_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_d_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_D_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_d_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_D_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_d_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_D_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_d_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.cpu_E_jtag_debug_module_address                       (mm_interconnect_0_cpu_e_jtag_debug_module_address),      //                         cpu_E_jtag_debug_module.address
		.cpu_E_jtag_debug_module_write                         (mm_interconnect_0_cpu_e_jtag_debug_module_write),        //                                                .write
		.cpu_E_jtag_debug_module_read                          (mm_interconnect_0_cpu_e_jtag_debug_module_read),         //                                                .read
		.cpu_E_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_e_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_E_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_e_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_E_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_e_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_E_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_e_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_E_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_e_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.cpu_F_jtag_debug_module_address                       (mm_interconnect_0_cpu_f_jtag_debug_module_address),      //                         cpu_F_jtag_debug_module.address
		.cpu_F_jtag_debug_module_write                         (mm_interconnect_0_cpu_f_jtag_debug_module_write),        //                                                .write
		.cpu_F_jtag_debug_module_read                          (mm_interconnect_0_cpu_f_jtag_debug_module_read),         //                                                .read
		.cpu_F_jtag_debug_module_readdata                      (mm_interconnect_0_cpu_f_jtag_debug_module_readdata),     //                                                .readdata
		.cpu_F_jtag_debug_module_writedata                     (mm_interconnect_0_cpu_f_jtag_debug_module_writedata),    //                                                .writedata
		.cpu_F_jtag_debug_module_byteenable                    (mm_interconnect_0_cpu_f_jtag_debug_module_byteenable),   //                                                .byteenable
		.cpu_F_jtag_debug_module_waitrequest                   (mm_interconnect_0_cpu_f_jtag_debug_module_waitrequest),  //                                                .waitrequest
		.cpu_F_jtag_debug_module_debugaccess                   (mm_interconnect_0_cpu_f_jtag_debug_module_debugaccess),  //                                                .debugaccess
		.fifo_AB_0_in_write                                    (mm_interconnect_0_fifo_ab_0_in_write),                   //                                    fifo_AB_0_in.write
		.fifo_AB_0_in_writedata                                (mm_interconnect_0_fifo_ab_0_in_writedata),               //                                                .writedata
		.fifo_AB_0_in_waitrequest                              (mm_interconnect_0_fifo_ab_0_in_waitrequest),             //                                                .waitrequest
		.fifo_AB_0_in_csr_address                              (mm_interconnect_0_fifo_ab_0_in_csr_address),             //                                fifo_AB_0_in_csr.address
		.fifo_AB_0_in_csr_write                                (mm_interconnect_0_fifo_ab_0_in_csr_write),               //                                                .write
		.fifo_AB_0_in_csr_read                                 (mm_interconnect_0_fifo_ab_0_in_csr_read),                //                                                .read
		.fifo_AB_0_in_csr_readdata                             (mm_interconnect_0_fifo_ab_0_in_csr_readdata),            //                                                .readdata
		.fifo_AB_0_in_csr_writedata                            (mm_interconnect_0_fifo_ab_0_in_csr_writedata),           //                                                .writedata
		.fifo_AB_0_out_read                                    (mm_interconnect_0_fifo_ab_0_out_read),                   //                                   fifo_AB_0_out.read
		.fifo_AB_0_out_readdata                                (mm_interconnect_0_fifo_ab_0_out_readdata),               //                                                .readdata
		.fifo_AB_0_out_waitrequest                             (mm_interconnect_0_fifo_ab_0_out_waitrequest),            //                                                .waitrequest
		.fifo_AB_1_in_write                                    (mm_interconnect_0_fifo_ab_1_in_write),                   //                                    fifo_AB_1_in.write
		.fifo_AB_1_in_writedata                                (mm_interconnect_0_fifo_ab_1_in_writedata),               //                                                .writedata
		.fifo_AB_1_in_waitrequest                              (mm_interconnect_0_fifo_ab_1_in_waitrequest),             //                                                .waitrequest
		.fifo_AB_1_in_csr_address                              (mm_interconnect_0_fifo_ab_1_in_csr_address),             //                                fifo_AB_1_in_csr.address
		.fifo_AB_1_in_csr_write                                (mm_interconnect_0_fifo_ab_1_in_csr_write),               //                                                .write
		.fifo_AB_1_in_csr_read                                 (mm_interconnect_0_fifo_ab_1_in_csr_read),                //                                                .read
		.fifo_AB_1_in_csr_readdata                             (mm_interconnect_0_fifo_ab_1_in_csr_readdata),            //                                                .readdata
		.fifo_AB_1_in_csr_writedata                            (mm_interconnect_0_fifo_ab_1_in_csr_writedata),           //                                                .writedata
		.fifo_AB_1_out_read                                    (mm_interconnect_0_fifo_ab_1_out_read),                   //                                   fifo_AB_1_out.read
		.fifo_AB_1_out_readdata                                (mm_interconnect_0_fifo_ab_1_out_readdata),               //                                                .readdata
		.fifo_AB_1_out_waitrequest                             (mm_interconnect_0_fifo_ab_1_out_waitrequest),            //                                                .waitrequest
		.fifo_AB_2_in_write                                    (mm_interconnect_0_fifo_ab_2_in_write),                   //                                    fifo_AB_2_in.write
		.fifo_AB_2_in_writedata                                (mm_interconnect_0_fifo_ab_2_in_writedata),               //                                                .writedata
		.fifo_AB_2_in_waitrequest                              (mm_interconnect_0_fifo_ab_2_in_waitrequest),             //                                                .waitrequest
		.fifo_AB_2_in_csr_address                              (mm_interconnect_0_fifo_ab_2_in_csr_address),             //                                fifo_AB_2_in_csr.address
		.fifo_AB_2_in_csr_write                                (mm_interconnect_0_fifo_ab_2_in_csr_write),               //                                                .write
		.fifo_AB_2_in_csr_read                                 (mm_interconnect_0_fifo_ab_2_in_csr_read),                //                                                .read
		.fifo_AB_2_in_csr_readdata                             (mm_interconnect_0_fifo_ab_2_in_csr_readdata),            //                                                .readdata
		.fifo_AB_2_in_csr_writedata                            (mm_interconnect_0_fifo_ab_2_in_csr_writedata),           //                                                .writedata
		.fifo_AB_2_out_read                                    (mm_interconnect_0_fifo_ab_2_out_read),                   //                                   fifo_AB_2_out.read
		.fifo_AB_2_out_readdata                                (mm_interconnect_0_fifo_ab_2_out_readdata),               //                                                .readdata
		.fifo_AB_2_out_waitrequest                             (mm_interconnect_0_fifo_ab_2_out_waitrequest),            //                                                .waitrequest
		.fifo_AD_in_write                                      (mm_interconnect_0_fifo_ad_in_write),                     //                                      fifo_AD_in.write
		.fifo_AD_in_writedata                                  (mm_interconnect_0_fifo_ad_in_writedata),                 //                                                .writedata
		.fifo_AD_in_waitrequest                                (mm_interconnect_0_fifo_ad_in_waitrequest),               //                                                .waitrequest
		.fifo_AD_in_csr_address                                (mm_interconnect_0_fifo_ad_in_csr_address),               //                                  fifo_AD_in_csr.address
		.fifo_AD_in_csr_write                                  (mm_interconnect_0_fifo_ad_in_csr_write),                 //                                                .write
		.fifo_AD_in_csr_read                                   (mm_interconnect_0_fifo_ad_in_csr_read),                  //                                                .read
		.fifo_AD_in_csr_readdata                               (mm_interconnect_0_fifo_ad_in_csr_readdata),              //                                                .readdata
		.fifo_AD_in_csr_writedata                              (mm_interconnect_0_fifo_ad_in_csr_writedata),             //                                                .writedata
		.fifo_AD_out_read                                      (mm_interconnect_0_fifo_ad_out_read),                     //                                     fifo_AD_out.read
		.fifo_AD_out_readdata                                  (mm_interconnect_0_fifo_ad_out_readdata),                 //                                                .readdata
		.fifo_AD_out_waitrequest                               (mm_interconnect_0_fifo_ad_out_waitrequest),              //                                                .waitrequest
		.fifo_AE_in_write                                      (mm_interconnect_0_fifo_ae_in_write),                     //                                      fifo_AE_in.write
		.fifo_AE_in_writedata                                  (mm_interconnect_0_fifo_ae_in_writedata),                 //                                                .writedata
		.fifo_AE_in_waitrequest                                (mm_interconnect_0_fifo_ae_in_waitrequest),               //                                                .waitrequest
		.fifo_AE_in_csr_address                                (mm_interconnect_0_fifo_ae_in_csr_address),               //                                  fifo_AE_in_csr.address
		.fifo_AE_in_csr_write                                  (mm_interconnect_0_fifo_ae_in_csr_write),                 //                                                .write
		.fifo_AE_in_csr_read                                   (mm_interconnect_0_fifo_ae_in_csr_read),                  //                                                .read
		.fifo_AE_in_csr_readdata                               (mm_interconnect_0_fifo_ae_in_csr_readdata),              //                                                .readdata
		.fifo_AE_in_csr_writedata                              (mm_interconnect_0_fifo_ae_in_csr_writedata),             //                                                .writedata
		.fifo_AE_out_read                                      (mm_interconnect_0_fifo_ae_out_read),                     //                                     fifo_AE_out.read
		.fifo_AE_out_readdata                                  (mm_interconnect_0_fifo_ae_out_readdata),                 //                                                .readdata
		.fifo_AE_out_waitrequest                               (mm_interconnect_0_fifo_ae_out_waitrequest),              //                                                .waitrequest
		.fifo_AF_in_write                                      (mm_interconnect_0_fifo_af_in_write),                     //                                      fifo_AF_in.write
		.fifo_AF_in_writedata                                  (mm_interconnect_0_fifo_af_in_writedata),                 //                                                .writedata
		.fifo_AF_in_waitrequest                                (mm_interconnect_0_fifo_af_in_waitrequest),               //                                                .waitrequest
		.fifo_AF_in_csr_address                                (mm_interconnect_0_fifo_af_in_csr_address),               //                                  fifo_AF_in_csr.address
		.fifo_AF_in_csr_write                                  (mm_interconnect_0_fifo_af_in_csr_write),                 //                                                .write
		.fifo_AF_in_csr_read                                   (mm_interconnect_0_fifo_af_in_csr_read),                  //                                                .read
		.fifo_AF_in_csr_readdata                               (mm_interconnect_0_fifo_af_in_csr_readdata),              //                                                .readdata
		.fifo_AF_in_csr_writedata                              (mm_interconnect_0_fifo_af_in_csr_writedata),             //                                                .writedata
		.fifo_AF_out_read                                      (mm_interconnect_0_fifo_af_out_read),                     //                                     fifo_AF_out.read
		.fifo_AF_out_readdata                                  (mm_interconnect_0_fifo_af_out_readdata),                 //                                                .readdata
		.fifo_AF_out_waitrequest                               (mm_interconnect_0_fifo_af_out_waitrequest),              //                                                .waitrequest
		.fifo_BC_in_write                                      (mm_interconnect_0_fifo_bc_in_write),                     //                                      fifo_BC_in.write
		.fifo_BC_in_writedata                                  (mm_interconnect_0_fifo_bc_in_writedata),                 //                                                .writedata
		.fifo_BC_in_waitrequest                                (mm_interconnect_0_fifo_bc_in_waitrequest),               //                                                .waitrequest
		.fifo_BC_in_csr_address                                (mm_interconnect_0_fifo_bc_in_csr_address),               //                                  fifo_BC_in_csr.address
		.fifo_BC_in_csr_write                                  (mm_interconnect_0_fifo_bc_in_csr_write),                 //                                                .write
		.fifo_BC_in_csr_read                                   (mm_interconnect_0_fifo_bc_in_csr_read),                  //                                                .read
		.fifo_BC_in_csr_readdata                               (mm_interconnect_0_fifo_bc_in_csr_readdata),              //                                                .readdata
		.fifo_BC_in_csr_writedata                              (mm_interconnect_0_fifo_bc_in_csr_writedata),             //                                                .writedata
		.fifo_BC_out_read                                      (mm_interconnect_0_fifo_bc_out_read),                     //                                     fifo_BC_out.read
		.fifo_BC_out_readdata                                  (mm_interconnect_0_fifo_bc_out_readdata),                 //                                                .readdata
		.fifo_BC_out_waitrequest                               (mm_interconnect_0_fifo_bc_out_waitrequest),              //                                                .waitrequest
		.fifo_CD_in_write                                      (mm_interconnect_0_fifo_cd_in_write),                     //                                      fifo_CD_in.write
		.fifo_CD_in_writedata                                  (mm_interconnect_0_fifo_cd_in_writedata),                 //                                                .writedata
		.fifo_CD_in_waitrequest                                (mm_interconnect_0_fifo_cd_in_waitrequest),               //                                                .waitrequest
		.fifo_CD_in_csr_address                                (mm_interconnect_0_fifo_cd_in_csr_address),               //                                  fifo_CD_in_csr.address
		.fifo_CD_in_csr_write                                  (mm_interconnect_0_fifo_cd_in_csr_write),                 //                                                .write
		.fifo_CD_in_csr_read                                   (mm_interconnect_0_fifo_cd_in_csr_read),                  //                                                .read
		.fifo_CD_in_csr_readdata                               (mm_interconnect_0_fifo_cd_in_csr_readdata),              //                                                .readdata
		.fifo_CD_in_csr_writedata                              (mm_interconnect_0_fifo_cd_in_csr_writedata),             //                                                .writedata
		.fifo_CD_out_read                                      (mm_interconnect_0_fifo_cd_out_read),                     //                                     fifo_CD_out.read
		.fifo_CD_out_readdata                                  (mm_interconnect_0_fifo_cd_out_readdata),                 //                                                .readdata
		.fifo_CD_out_waitrequest                               (mm_interconnect_0_fifo_cd_out_waitrequest),              //                                                .waitrequest
		.fifo_DE_in_write                                      (mm_interconnect_0_fifo_de_in_write),                     //                                      fifo_DE_in.write
		.fifo_DE_in_writedata                                  (mm_interconnect_0_fifo_de_in_writedata),                 //                                                .writedata
		.fifo_DE_in_waitrequest                                (mm_interconnect_0_fifo_de_in_waitrequest),               //                                                .waitrequest
		.fifo_DE_in_csr_address                                (mm_interconnect_0_fifo_de_in_csr_address),               //                                  fifo_DE_in_csr.address
		.fifo_DE_in_csr_write                                  (mm_interconnect_0_fifo_de_in_csr_write),                 //                                                .write
		.fifo_DE_in_csr_read                                   (mm_interconnect_0_fifo_de_in_csr_read),                  //                                                .read
		.fifo_DE_in_csr_readdata                               (mm_interconnect_0_fifo_de_in_csr_readdata),              //                                                .readdata
		.fifo_DE_in_csr_writedata                              (mm_interconnect_0_fifo_de_in_csr_writedata),             //                                                .writedata
		.fifo_DE_out_read                                      (mm_interconnect_0_fifo_de_out_read),                     //                                     fifo_DE_out.read
		.fifo_DE_out_readdata                                  (mm_interconnect_0_fifo_de_out_readdata),                 //                                                .readdata
		.fifo_DE_out_waitrequest                               (mm_interconnect_0_fifo_de_out_waitrequest),              //                                                .waitrequest
		.fifo_EF_in_write                                      (mm_interconnect_0_fifo_ef_in_write),                     //                                      fifo_EF_in.write
		.fifo_EF_in_writedata                                  (mm_interconnect_0_fifo_ef_in_writedata),                 //                                                .writedata
		.fifo_EF_in_waitrequest                                (mm_interconnect_0_fifo_ef_in_waitrequest),               //                                                .waitrequest
		.fifo_EF_in_csr_address                                (mm_interconnect_0_fifo_ef_in_csr_address),               //                                  fifo_EF_in_csr.address
		.fifo_EF_in_csr_write                                  (mm_interconnect_0_fifo_ef_in_csr_write),                 //                                                .write
		.fifo_EF_in_csr_read                                   (mm_interconnect_0_fifo_ef_in_csr_read),                  //                                                .read
		.fifo_EF_in_csr_readdata                               (mm_interconnect_0_fifo_ef_in_csr_readdata),              //                                                .readdata
		.fifo_EF_in_csr_writedata                              (mm_interconnect_0_fifo_ef_in_csr_writedata),             //                                                .writedata
		.fifo_EF_out_read                                      (mm_interconnect_0_fifo_ef_out_read),                     //                                     fifo_EF_out.read
		.fifo_EF_out_readdata                                  (mm_interconnect_0_fifo_ef_out_readdata),                 //                                                .readdata
		.fifo_EF_out_waitrequest                               (mm_interconnect_0_fifo_ef_out_waitrequest),              //                                                .waitrequest
		.highTimer_A_s1_address                                (mm_interconnect_0_hightimer_a_s1_address),               //                                  highTimer_A_s1.address
		.highTimer_A_s1_write                                  (mm_interconnect_0_hightimer_a_s1_write),                 //                                                .write
		.highTimer_A_s1_readdata                               (mm_interconnect_0_hightimer_a_s1_readdata),              //                                                .readdata
		.highTimer_A_s1_writedata                              (mm_interconnect_0_hightimer_a_s1_writedata),             //                                                .writedata
		.highTimer_A_s1_chipselect                             (mm_interconnect_0_hightimer_a_s1_chipselect),            //                                                .chipselect
		.highTimer_B_s1_address                                (mm_interconnect_0_hightimer_b_s1_address),               //                                  highTimer_B_s1.address
		.highTimer_B_s1_write                                  (mm_interconnect_0_hightimer_b_s1_write),                 //                                                .write
		.highTimer_B_s1_readdata                               (mm_interconnect_0_hightimer_b_s1_readdata),              //                                                .readdata
		.highTimer_B_s1_writedata                              (mm_interconnect_0_hightimer_b_s1_writedata),             //                                                .writedata
		.highTimer_B_s1_chipselect                             (mm_interconnect_0_hightimer_b_s1_chipselect),            //                                                .chipselect
		.highTimer_C_s1_address                                (mm_interconnect_0_hightimer_c_s1_address),               //                                  highTimer_C_s1.address
		.highTimer_C_s1_write                                  (mm_interconnect_0_hightimer_c_s1_write),                 //                                                .write
		.highTimer_C_s1_readdata                               (mm_interconnect_0_hightimer_c_s1_readdata),              //                                                .readdata
		.highTimer_C_s1_writedata                              (mm_interconnect_0_hightimer_c_s1_writedata),             //                                                .writedata
		.highTimer_C_s1_chipselect                             (mm_interconnect_0_hightimer_c_s1_chipselect),            //                                                .chipselect
		.highTimer_D_s1_address                                (mm_interconnect_0_hightimer_d_s1_address),               //                                  highTimer_D_s1.address
		.highTimer_D_s1_write                                  (mm_interconnect_0_hightimer_d_s1_write),                 //                                                .write
		.highTimer_D_s1_readdata                               (mm_interconnect_0_hightimer_d_s1_readdata),              //                                                .readdata
		.highTimer_D_s1_writedata                              (mm_interconnect_0_hightimer_d_s1_writedata),             //                                                .writedata
		.highTimer_D_s1_chipselect                             (mm_interconnect_0_hightimer_d_s1_chipselect),            //                                                .chipselect
		.highTimer_E_s1_address                                (mm_interconnect_0_hightimer_e_s1_address),               //                                  highTimer_E_s1.address
		.highTimer_E_s1_write                                  (mm_interconnect_0_hightimer_e_s1_write),                 //                                                .write
		.highTimer_E_s1_readdata                               (mm_interconnect_0_hightimer_e_s1_readdata),              //                                                .readdata
		.highTimer_E_s1_writedata                              (mm_interconnect_0_hightimer_e_s1_writedata),             //                                                .writedata
		.highTimer_E_s1_chipselect                             (mm_interconnect_0_hightimer_e_s1_chipselect),            //                                                .chipselect
		.highTimer_F_s1_address                                (mm_interconnect_0_hightimer_f_s1_address),               //                                  highTimer_F_s1.address
		.highTimer_F_s1_write                                  (mm_interconnect_0_hightimer_f_s1_write),                 //                                                .write
		.highTimer_F_s1_readdata                               (mm_interconnect_0_hightimer_f_s1_readdata),              //                                                .readdata
		.highTimer_F_s1_writedata                              (mm_interconnect_0_hightimer_f_s1_writedata),             //                                                .writedata
		.highTimer_F_s1_chipselect                             (mm_interconnect_0_hightimer_f_s1_chipselect),            //                                                .chipselect
		.jtag_A_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_a_avalon_jtag_slave_address),     //                        jtag_A_avalon_jtag_slave.address
		.jtag_A_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_a_avalon_jtag_slave_write),       //                                                .write
		.jtag_A_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_a_avalon_jtag_slave_read),        //                                                .read
		.jtag_A_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_a_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_A_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_a_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_A_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_a_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_A_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_a_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_B_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_b_avalon_jtag_slave_address),     //                        jtag_B_avalon_jtag_slave.address
		.jtag_B_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_b_avalon_jtag_slave_write),       //                                                .write
		.jtag_B_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_b_avalon_jtag_slave_read),        //                                                .read
		.jtag_B_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_b_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_B_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_b_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_B_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_b_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_B_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_b_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_C_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_c_avalon_jtag_slave_address),     //                        jtag_C_avalon_jtag_slave.address
		.jtag_C_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_c_avalon_jtag_slave_write),       //                                                .write
		.jtag_C_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_c_avalon_jtag_slave_read),        //                                                .read
		.jtag_C_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_c_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_C_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_c_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_C_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_c_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_C_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_c_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_D_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_d_avalon_jtag_slave_address),     //                        jtag_D_avalon_jtag_slave.address
		.jtag_D_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_d_avalon_jtag_slave_write),       //                                                .write
		.jtag_D_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_d_avalon_jtag_slave_read),        //                                                .read
		.jtag_D_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_d_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_D_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_d_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_D_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_d_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_D_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_d_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_E_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_e_avalon_jtag_slave_address),     //                        jtag_E_avalon_jtag_slave.address
		.jtag_E_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_e_avalon_jtag_slave_write),       //                                                .write
		.jtag_E_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_e_avalon_jtag_slave_read),        //                                                .read
		.jtag_E_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_e_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_E_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_e_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_E_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_e_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_E_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_e_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_F_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_f_avalon_jtag_slave_address),     //                        jtag_F_avalon_jtag_slave.address
		.jtag_F_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_f_avalon_jtag_slave_write),       //                                                .write
		.jtag_F_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_f_avalon_jtag_slave_read),        //                                                .read
		.jtag_F_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_f_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_F_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_f_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_F_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_f_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_F_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_f_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.led_out_s1_address                                    (mm_interconnect_0_led_out_s1_address),                   //                                      led_out_s1.address
		.led_out_s1_write                                      (mm_interconnect_0_led_out_s1_write),                     //                                                .write
		.led_out_s1_readdata                                   (mm_interconnect_0_led_out_s1_readdata),                  //                                                .readdata
		.led_out_s1_writedata                                  (mm_interconnect_0_led_out_s1_writedata),                 //                                                .writedata
		.led_out_s1_chipselect                                 (mm_interconnect_0_led_out_s1_chipselect),                //                                                .chipselect
		.PLL_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                //                                   PLL_pll_slave.address
		.PLL_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                  //                                                .write
		.PLL_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                   //                                                .read
		.PLL_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),               //                                                .readdata
		.PLL_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),              //                                                .writedata
		.SDRAM_controller_s1_address                           (mm_interconnect_0_sdram_controller_s1_address),          //                             SDRAM_controller_s1.address
		.SDRAM_controller_s1_write                             (mm_interconnect_0_sdram_controller_s1_write),            //                                                .write
		.SDRAM_controller_s1_read                              (mm_interconnect_0_sdram_controller_s1_read),             //                                                .read
		.SDRAM_controller_s1_readdata                          (mm_interconnect_0_sdram_controller_s1_readdata),         //                                                .readdata
		.SDRAM_controller_s1_writedata                         (mm_interconnect_0_sdram_controller_s1_writedata),        //                                                .writedata
		.SDRAM_controller_s1_byteenable                        (mm_interconnect_0_sdram_controller_s1_byteenable),       //                                                .byteenable
		.SDRAM_controller_s1_readdatavalid                     (mm_interconnect_0_sdram_controller_s1_readdatavalid),    //                                                .readdatavalid
		.SDRAM_controller_s1_waitrequest                       (mm_interconnect_0_sdram_controller_s1_waitrequest),      //                                                .waitrequest
		.SDRAM_controller_s1_chipselect                        (mm_interconnect_0_sdram_controller_s1_chipselect),       //                                                .chipselect
		.sysid_A_control_slave_address                         (mm_interconnect_0_sysid_a_control_slave_address),        //                           sysid_A_control_slave.address
		.sysid_A_control_slave_readdata                        (mm_interconnect_0_sysid_a_control_slave_readdata),       //                                                .readdata
		.sysid_B_control_slave_address                         (mm_interconnect_0_sysid_b_control_slave_address),        //                           sysid_B_control_slave.address
		.sysid_B_control_slave_readdata                        (mm_interconnect_0_sysid_b_control_slave_readdata),       //                                                .readdata
		.sysid_C_control_slave_address                         (mm_interconnect_0_sysid_c_control_slave_address),        //                           sysid_C_control_slave.address
		.sysid_C_control_slave_readdata                        (mm_interconnect_0_sysid_c_control_slave_readdata),       //                                                .readdata
		.sysid_D_control_slave_address                         (mm_interconnect_0_sysid_d_control_slave_address),        //                           sysid_D_control_slave.address
		.sysid_D_control_slave_readdata                        (mm_interconnect_0_sysid_d_control_slave_readdata),       //                                                .readdata
		.sysid_E_control_slave_address                         (mm_interconnect_0_sysid_e_control_slave_address),        //                           sysid_E_control_slave.address
		.sysid_E_control_slave_readdata                        (mm_interconnect_0_sysid_e_control_slave_readdata),       //                                                .readdata
		.sysid_F_control_slave_address                         (mm_interconnect_0_sysid_f_control_slave_address),        //                           sysid_F_control_slave.address
		.sysid_F_control_slave_readdata                        (mm_interconnect_0_sysid_f_control_slave_readdata),       //                                                .readdata
		.timer_A_s1_address                                    (mm_interconnect_0_timer_a_s1_address),                   //                                      timer_A_s1.address
		.timer_A_s1_write                                      (mm_interconnect_0_timer_a_s1_write),                     //                                                .write
		.timer_A_s1_readdata                                   (mm_interconnect_0_timer_a_s1_readdata),                  //                                                .readdata
		.timer_A_s1_writedata                                  (mm_interconnect_0_timer_a_s1_writedata),                 //                                                .writedata
		.timer_A_s1_chipselect                                 (mm_interconnect_0_timer_a_s1_chipselect),                //                                                .chipselect
		.timer_B_s1_address                                    (mm_interconnect_0_timer_b_s1_address),                   //                                      timer_B_s1.address
		.timer_B_s1_write                                      (mm_interconnect_0_timer_b_s1_write),                     //                                                .write
		.timer_B_s1_readdata                                   (mm_interconnect_0_timer_b_s1_readdata),                  //                                                .readdata
		.timer_B_s1_writedata                                  (mm_interconnect_0_timer_b_s1_writedata),                 //                                                .writedata
		.timer_B_s1_chipselect                                 (mm_interconnect_0_timer_b_s1_chipselect),                //                                                .chipselect
		.timer_C_s1_address                                    (mm_interconnect_0_timer_c_s1_address),                   //                                      timer_C_s1.address
		.timer_C_s1_write                                      (mm_interconnect_0_timer_c_s1_write),                     //                                                .write
		.timer_C_s1_readdata                                   (mm_interconnect_0_timer_c_s1_readdata),                  //                                                .readdata
		.timer_C_s1_writedata                                  (mm_interconnect_0_timer_c_s1_writedata),                 //                                                .writedata
		.timer_C_s1_chipselect                                 (mm_interconnect_0_timer_c_s1_chipselect),                //                                                .chipselect
		.timer_D_s1_address                                    (mm_interconnect_0_timer_d_s1_address),                   //                                      timer_D_s1.address
		.timer_D_s1_write                                      (mm_interconnect_0_timer_d_s1_write),                     //                                                .write
		.timer_D_s1_readdata                                   (mm_interconnect_0_timer_d_s1_readdata),                  //                                                .readdata
		.timer_D_s1_writedata                                  (mm_interconnect_0_timer_d_s1_writedata),                 //                                                .writedata
		.timer_D_s1_chipselect                                 (mm_interconnect_0_timer_d_s1_chipselect),                //                                                .chipselect
		.timer_E_s1_address                                    (mm_interconnect_0_timer_e_s1_address),                   //                                      timer_E_s1.address
		.timer_E_s1_write                                      (mm_interconnect_0_timer_e_s1_write),                     //                                                .write
		.timer_E_s1_readdata                                   (mm_interconnect_0_timer_e_s1_readdata),                  //                                                .readdata
		.timer_E_s1_writedata                                  (mm_interconnect_0_timer_e_s1_writedata),                 //                                                .writedata
		.timer_E_s1_chipselect                                 (mm_interconnect_0_timer_e_s1_chipselect),                //                                                .chipselect
		.timer_F_s1_address                                    (mm_interconnect_0_timer_f_s1_address),                   //                                      timer_F_s1.address
		.timer_F_s1_write                                      (mm_interconnect_0_timer_f_s1_write),                     //                                                .write
		.timer_F_s1_readdata                                   (mm_interconnect_0_timer_f_s1_readdata),                  //                                                .readdata
		.timer_F_s1_writedata                                  (mm_interconnect_0_timer_f_s1_writedata),                 //                                                .writedata
		.timer_F_s1_chipselect                                 (mm_interconnect_0_timer_f_s1_chipselect)                 //                                                .chipselect
	);

	HwJSoC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),           // receiver8.irq
		.sender_irq    (cpu_a_d_irq_irq)                     //    sender.irq
	);

	HwJSoC_irq_mapper_001 irq_mapper_001 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_b_d_irq_irq)                     //    sender.irq
	);

	HwJSoC_irq_mapper_001 irq_mapper_002 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_005_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_002_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_002_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_c_d_irq_irq)                     //    sender.irq
	);

	HwJSoC_irq_mapper_003 irq_mapper_003 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_006_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_003_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_003_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver6_irq),           // receiver4.irq
		.sender_irq    (cpu_d_d_irq_irq)                     //    sender.irq
	);

	HwJSoC_irq_mapper_001 irq_mapper_004 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_007_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_004_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_004_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_e_d_irq_irq)                     //    sender.irq
	);

	HwJSoC_irq_mapper_005 irq_mapper_005 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_008_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_005_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_005_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_005_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_f_d_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (7),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_a_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_c_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3      (cpu_d_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4      (cpu_b_jtag_debug_module_reset_reset), // reset_in4.reset
		.reset_in5      (cpu_e_jtag_debug_module_reset_reset), // reset_in5.reset
		.reset_in6      (cpu_f_jtag_debug_module_reset_reset), // reset_in6.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_a_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_a_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_b_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_b_jtag_debug_module_reset_reset),    // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (cpu_c_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_005_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (cpu_d_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_006_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (cpu_e_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_007_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (cpu_f_jtag_debug_module_reset_reset),    // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_008_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_a_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_d_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_010 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_a_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_e_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_010_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_011 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_a_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_f_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_011_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_012 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_b_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_c_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_012_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_013 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_c_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_d_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_013_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_014 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_d_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_e_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_014_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_015 (
		.reset_in0      (cpu_e_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                      // reset_in1.reset
		.reset_in2      (cpu_f_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_015_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
